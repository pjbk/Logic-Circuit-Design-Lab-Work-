CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
14 Logic Display~
6 791 125 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
43809.8 14
0
8 2-In OR~
219 628 143 0 3 22
0 13 12 11
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
842 0 0
2
43809.8 13
0
10 2-In NAND~
219 697 272 0 3 22
0 9 10 8
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3277 0 0
2
43809.8 12
0
10 2-In NAND~
219 612 319 0 3 22
0 6 6 10
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4212 0 0
2
43809.8 11
0
10 2-In NAND~
219 607 241 0 3 22
0 7 7 9
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4720 0 0
2
43809.8 10
0
14 Logic Display~
6 797 249 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5551 0 0
2
43809.8 9
0
9 2-In NOR~
219 612 420 0 3 22
0 5 4 2
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6986 0 0
2
43809.8 8
0
9 2-In NOR~
219 717 420 0 3 22
0 2 2 3
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8745 0 0
2
43809.8 7
0
14 Logic Display~
6 806 402 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
43809.8 6
0
13 Logic Switch~
5 490 119 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
43809.8 5
0
13 Logic Switch~
5 491 167 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
43809.8 4
0
13 Logic Switch~
5 496 232 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
631 0 0
2
43809.8 3
0
13 Logic Switch~
5 498 328 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9466 0 0
2
43809.8 2
0
13 Logic Switch~
5 507 397 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3266 0 0
2
43809.8 1
0
13 Logic Switch~
5 505 442 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
43809.8 0
0
15
0 2 2 0 0 16 0 0 8 3 0 3
666 420
666 429
704 429
3 1 3 0 0 16 0 8 9 0 0 2
756 420
806 420
3 1 2 0 0 16 0 7 8 0 0 4
651 420
666 420
666 411
704 411
1 2 4 0 0 16 0 15 7 0 0 4
517 442
589 442
589 429
599 429
1 1 5 0 0 16 0 14 7 0 0 4
519 397
589 397
589 411
599 411
0 1 6 0 0 16 0 0 4 11 0 3
564 328
564 310
588 310
0 2 7 0 0 16 0 0 5 12 0 3
545 232
545 250
583 250
3 1 8 0 0 16 0 3 6 0 0 3
724 272
797 272
797 267
3 1 9 0 0 16 0 5 3 0 0 4
634 241
665 241
665 263
673 263
3 2 10 0 0 16 0 4 3 0 0 4
639 319
665 319
665 281
673 281
1 2 6 0 0 16 0 13 4 0 0 2
510 328
588 328
1 1 7 0 0 16 0 12 5 0 0 2
508 232
583 232
3 1 11 0 0 16 0 2 1 0 0 2
661 143
791 143
1 2 12 0 0 16 0 11 2 0 0 4
503 167
579 167
579 152
615 152
1 1 13 0 0 16 0 10 2 0 0 4
502 119
579 119
579 134
615 134
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
299 124 424 148
309 131 413 147
13 Basic OR gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
262 263 507 287
272 271 496 287
28 OR gate using Universal NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
256 405 493 429
266 413 482 429
27 OR gate using Universal NOR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
