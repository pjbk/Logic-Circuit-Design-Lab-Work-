CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 102 552 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
43557.5 0
0
13 Logic Switch~
5 101 478 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
43557.5 1
0
13 Logic Switch~
5 103 420 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
43557.5 2
0
13 Logic Switch~
5 102 343 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3178 0 0
2
43557.5 3
0
13 Logic Switch~
5 101 303 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
43557.5 4
0
13 Logic Switch~
5 99 263 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
43557.5 5
0
13 Logic Switch~
5 101 224 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
43557.5 6
0
13 Logic Switch~
5 100 187 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
43557.5 7
0
13 Logic Switch~
5 100 151 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
43557.5 8
0
13 Logic Switch~
5 102 114 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
43557.5 9
0
13 Logic Switch~
5 101 65 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
43557.5 10
0
14 Logic Display~
6 1092 210 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
43557.5 11
0
5 4071~
219 968 232 0 3 22
0 18 17 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
9281 0 0
2
43557.5 12
0
8 4-In OR~
219 850 220 0 5 22
0 22 21 20 19 18
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
8464 0 0
2
43557.5 13
0
8 4-In OR~
219 697 205 0 5 22
0 26 25 24 23 22
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
7168 0 0
2
43557.5 14
0
5 4082~
219 365 413 0 5 22
0 3 11 13 12 17
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3171 0 0
2
43557.5 15
0
5 4082~
219 365 363 0 5 22
0 4 11 13 14 19
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
4139 0 0
2
43557.5 16
0
5 4082~
219 365 313 0 5 22
0 5 11 15 12 20
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
6435 0 0
2
43557.5 17
0
5 4082~
219 361 264 0 5 22
0 6 11 15 14 21
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
5283 0 0
2
43557.5 18
0
5 4082~
219 362 205 0 5 22
0 7 16 12 13 23
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
6874 0 0
2
43557.5 19
0
5 4082~
219 361 152 0 5 22
0 8 16 13 14 24
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
5305 0 0
2
43557.5 20
0
5 4082~
219 363 98 0 5 22
0 9 16 15 12 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
34 0 0
2
43557.5 21
0
5 4082~
219 360 45 0 5 22
0 10 16 15 14 26
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
969 0 0
2
43557.5 22
0
5 4049~
219 204 548 0 2 22
0 12 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
8402 0 0
2
43557.5 23
0
5 4049~
219 203 485 0 2 22
0 13 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3751 0 0
2
43557.5 24
0
5 4049~
219 206 425 0 2 22
0 11 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4292 0 0
2
43557.5 25
0
46
3 1 2 0 0 4224 0 13 12 0 0 3
1001 232
1092 232
1092 228
1 1 3 0 0 8320 0 4 16 0 0 5
114 343
114 390
328 390
328 400
341 400
1 1 4 0 0 8320 0 5 17 0 0 5
113 303
113 336
333 336
333 350
341 350
1 1 5 0 0 8320 0 6 18 0 0 5
111 263
111 289
333 289
333 300
341 300
1 1 6 0 0 8320 0 7 19 0 0 3
113 224
113 251
337 251
1 1 7 0 0 4224 0 8 20 0 0 4
112 187
330 187
330 192
338 192
1 1 8 0 0 8320 0 9 21 0 0 3
112 151
112 139
337 139
1 1 9 0 0 8320 0 10 22 0 0 3
114 114
114 85
339 85
1 1 10 0 0 8320 0 11 23 0 0 3
113 65
113 32
336 32
2 0 11 0 0 8320 0 16 0 0 21 3
341 409
341 408
131 408
0 4 12 0 0 4096 0 0 16 28 0 3
158 455
341 455
341 427
0 3 13 0 0 4096 0 0 16 27 0 4
149 438
333 438
333 418
341 418
0 4 14 0 0 4096 0 0 17 31 0 2
318 377
341 377
0 3 13 0 0 4096 0 0 17 27 0 2
149 368
341 368
0 2 11 0 0 0 0 0 17 21 0 2
131 359
341 359
0 4 12 0 0 0 0 0 18 28 0 2
158 327
341 327
0 3 15 0 0 4096 0 0 18 32 0 2
273 318
341 318
0 2 11 0 0 0 0 0 18 21 0 2
131 309
341 309
0 3 15 0 0 0 0 0 19 32 0 2
273 269
337 269
0 4 14 0 0 0 0 0 19 31 0 4
318 279
329 279
329 278
337 278
2 0 11 0 0 0 0 19 0 0 36 3
337 260
131 260
131 420
0 4 13 0 0 0 0 0 20 27 0 2
149 219
338 219
0 3 12 0 0 0 0 0 20 28 0 2
158 210
338 210
0 2 16 0 0 4096 0 0 20 33 0 2
238 201
338 201
0 2 16 0 0 0 0 0 21 33 0 4
238 149
329 149
329 148
337 148
0 4 14 0 0 0 0 0 21 31 0 2
318 166
337 166
0 3 13 0 0 4224 0 0 21 35 0 3
149 478
149 157
337 157
0 4 12 0 0 4224 0 0 22 34 0 3
158 552
158 112
339 112
0 3 15 0 0 0 0 0 22 32 0 2
273 103
339 103
0 2 16 0 0 4096 0 0 22 33 0 2
238 94
339 94
2 4 14 0 0 8320 0 24 23 0 0 4
225 548
318 548
318 59
336 59
2 3 15 0 0 8320 0 25 23 0 0 4
224 485
273 485
273 50
336 50
2 2 16 0 0 8320 0 26 23 0 0 4
227 425
238 425
238 41
336 41
1 1 12 0 0 0 0 1 24 0 0 4
114 552
181 552
181 548
189 548
1 1 13 0 0 0 0 2 25 0 0 4
113 478
180 478
180 485
188 485
1 1 11 0 0 0 0 3 26 0 0 4
115 420
183 420
183 425
191 425
5 2 17 0 0 4224 0 16 13 0 0 4
386 413
947 413
947 241
955 241
5 1 18 0 0 4224 0 14 13 0 0 4
883 220
948 220
948 223
955 223
4 5 19 0 0 4224 0 14 17 0 0 4
833 234
394 234
394 363
386 363
5 3 20 0 0 4224 0 18 14 0 0 4
386 313
820 313
820 225
833 225
5 2 21 0 0 4224 0 19 14 0 0 4
382 264
825 264
825 216
833 216
5 1 22 0 0 4224 0 15 14 0 0 4
730 205
825 205
825 207
833 207
5 4 23 0 0 4224 0 20 15 0 0 4
383 205
672 205
672 219
680 219
5 3 24 0 0 4224 0 21 15 0 0 4
382 152
662 152
662 210
680 210
5 2 25 0 0 4224 0 22 15 0 0 4
384 98
667 98
667 201
680 201
5 1 26 0 0 4224 0 23 15 0 0 4
381 45
672 45
672 192
680 192
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 175 71 199
44 183 60 199
2 I3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 214 87 238
60 222 76 238
2 I4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
29 147 66 171
39 155 55 171
2 I2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
27 99 64 123
37 107 53 123
2 I1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 257 87 281
60 265 76 281
2 I5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
46 289 83 313
56 297 72 313
2 I6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
43 335 80 359
53 343 69 359
2 I7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 52 73 76
46 60 62 76
2 I0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
42 408 79 432
52 416 68 432
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 460 75 484
48 468 64 484
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
33 530 70 554
43 538 59 554
2 S0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
