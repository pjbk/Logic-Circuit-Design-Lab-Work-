CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 309 281 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-53 -10 -46 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9395 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 309 385 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 C
-50 -18 -43 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3303 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 309 212 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-52 -7 -45 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4498 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 895 346 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9728 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 886 249 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 883 170 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3978 0 0
2
5.89774e-315 0
0
6 74136~
219 753 370 0 3 22
0 3 7 2
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3494 0 0
2
5.89774e-315 0
0
6 74136~
219 511 381 0 3 22
0 6 5 7
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3507 0 0
2
5.89774e-315 0
0
6 74136~
219 506 279 0 3 22
0 3 6 4
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5151 0 0
2
5.89774e-315 0
0
9
1 3 2 0 0 8320 0 4 7 0 0 3
895 364
895 370
786 370
1 0 3 0 0 8192 0 7 0 0 4 3
737 361
659 361
659 207
1 3 4 0 0 8320 0 5 9 0 0 3
886 267
886 279
539 279
1 0 3 0 0 8320 0 6 0 0 8 4
883 188
883 207
420 207
420 212
1 2 5 0 0 4224 0 2 8 0 0 4
321 385
487 385
487 390
495 390
1 1 6 0 0 4224 0 8 1 0 0 4
495 372
330 372
330 281
321 281
1 2 6 0 0 0 0 1 9 0 0 4
321 281
482 281
482 288
490 288
1 1 3 0 0 0 0 3 9 0 0 4
321 212
482 212
482 270
490 270
3 2 7 0 0 4224 0 8 7 0 0 4
544 381
729 381
729 379
737 379
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
832 338 861 362
842 346 850 362
1 z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
825 252 854 276
835 260 843 276
1 y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
822 178 851 202
832 186 840 202
1 x
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
