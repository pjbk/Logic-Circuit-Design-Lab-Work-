CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 313 334 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-59 -11 -38 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
42666.8 0
0
13 Logic Switch~
5 300 259 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-39 -8 -32 0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
42666.8 1
0
13 Logic Switch~
5 293 173 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-40 -8 -33 0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3221 0 0
2
42666.8 2
0
14 Logic Display~
6 1025 236 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
42666.8 3
0
14 Logic Display~
6 1022 159 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
42666.8 4
0
8 2-In OR~
219 914 254 0 3 22
0 4 5 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 Cout
59 -17 87 -9
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7121 0 0
2
42666.8 5
0
9 2-In AND~
219 740 246 0 3 22
0 7 6 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4484 0 0
2
42666.8 6
0
9 2-In AND~
219 565 246 0 3 22
0 9 8 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5996 0 0
2
42666.8 7
0
6 74136~
219 662 177 0 3 22
0 7 6 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 sum
306 -14 327 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7804 0 0
2
42666.8 8
0
6 74136~
219 446 173 0 3 22
0 9 8 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5523 0 0
2
42666.8 9
0
12
3 1 2 0 0 4224 0 6 4 0 0 2
947 254
1025 254
3 1 3 0 0 4224 0 9 5 0 0 2
695 177
1022 177
3 1 4 0 0 4224 0 7 6 0 0 4
761 246
893 246
893 245
901 245
3 2 5 0 0 12416 0 8 6 0 0 6
586 246
712 246
712 266
893 266
893 263
901 263
0 2 6 0 0 4096 0 0 7 9 0 2
638 255
716 255
0 1 7 0 0 8192 0 0 7 10 0 5
580 173
580 227
708 227
708 237
716 237
0 2 8 0 0 4224 0 0 8 11 0 2
422 255
541 255
0 1 9 0 0 8320 0 0 8 12 0 3
364 173
364 237
541 237
1 2 6 0 0 4224 0 1 9 0 0 4
325 334
638 334
638 186
646 186
3 1 7 0 0 4224 0 10 9 0 0 4
479 173
638 173
638 168
646 168
1 2 8 0 0 0 0 2 10 0 0 4
312 259
422 259
422 182
430 182
1 1 9 0 0 0 0 3 10 0 0 4
305 173
422 173
422 164
430 164
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
