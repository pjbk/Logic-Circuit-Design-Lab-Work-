CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 305 167 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3679 0 0
2
43550 5
0
13 Logic Switch~
5 316 237 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9342 0 0
2
43550 4
0
13 Logic Switch~
5 321 304 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3623 0 0
2
43550 3
0
13 Logic Switch~
5 374 469 0 1 11
0 4
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3722 0 0
2
43550 1
0
13 Logic Switch~
5 443 468 0 1 11
0 6
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8993 0 0
2
43550 0
0
9 Inverter~
13 353 321 0 2 22
0 3 2
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3723 0 0
2
43550 0
0
5 7415~
219 562 151 0 4 22
0 10 8 7 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
6244 0 0
2
43550 13
0
5 7415~
219 568 225 0 4 22
0 9 8 6 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
6421 0 0
2
43550 12
0
5 7415~
219 571 295 0 4 22
0 3 7 4 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
7743 0 0
2
43550 11
0
5 7415~
219 576 379 0 4 22
0 2 4 6 11
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
9840 0 0
2
43550 10
0
8 4-In OR~
219 746 251 0 5 22
0 14 13 12 11 5
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
6910 0 0
2
43550 9
0
9 Inverter~
13 372 424 0 2 22
0 4 8
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
449 0 0
2
43550 8
0
9 Inverter~
13 441 419 0 2 22
0 6 7
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8761 0 0
2
43550 7
0
14 Logic Display~
6 852 238 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6748 0 0
2
43550 6
0
20
2 1 2 0 0 8320 0 6 10 0 0 3
356 339
356 370
552 370
1 0 3 0 0 4096 0 6 0 0 10 2
356 303
356 304
0 3 4 0 0 4112 0 0 9 4 0 3
526 446
526 304
547 304
1 2 4 0 0 8336 0 12 10 0 0 5
375 442
375 446
539 446
539 379
552 379
5 1 5 0 0 4240 0 11 14 0 0 5
779 251
840 251
840 264
852 264
852 256
0 3 6 0 0 4240 0 0 8 7 0 3
503 441
503 234
544 234
1 3 6 0 0 16 0 13 10 0 0 5
444 437
444 441
544 441
544 388
552 388
0 2 7 0 0 4112 0 0 9 12 0 4
444 296
534 296
534 295
547 295
0 2 8 0 0 4112 0 0 8 13 0 2
375 225
544 225
1 1 3 0 0 4240 0 3 9 0 0 4
333 304
539 304
539 286
547 286
1 1 9 0 0 4240 0 2 8 0 0 4
328 237
536 237
536 216
544 216
2 3 7 0 0 4240 0 13 7 0 0 3
444 401
444 160
538 160
2 2 8 0 0 4240 0 12 7 0 0 3
375 406
375 151
538 151
1 1 10 0 0 4240 0 1 7 0 0 4
317 167
530 167
530 142
538 142
4 4 11 0 0 4240 0 10 11 0 0 4
597 379
716 379
716 265
729 265
4 3 12 0 0 4240 0 9 11 0 0 4
592 295
721 295
721 256
729 256
4 2 13 0 0 4240 0 8 11 0 0 4
589 225
716 225
716 247
729 247
4 1 14 0 0 4240 0 7 11 0 0 4
583 151
721 151
721 238
729 238
1 1 6 0 0 16 0 13 5 0 0 2
444 437
444 455
1 1 4 0 0 16 0 12 4 0 0 4
375 442
375 457
375 457
375 456
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
556 362 593 386
566 370 582 386
2 I3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
552 271 589 295
562 279 578 295
2 I2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
551 212 588 236
561 220 577 236
2 I1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
539 135 576 159
549 143 565 159
2 I0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
588 445 769 469
598 453 758 469
20 I0=0;I1=1;I2=A;I3=A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
334 501 523 525
344 509 512 525
21 F(A,B,C)=sum(1,3,5,6)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
