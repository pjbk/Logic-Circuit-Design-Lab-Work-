CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 243 220 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6901 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 240 155 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
842 0 0
2
5.89886e-315 0
0
9 Inverter~
13 987 224 0 2 22
0 5 2
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3277 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 737 100 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 775 98 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 811 99 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 845 98 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.89886e-315 0
0
5 7422~
219 944 287 0 5 22
0 4 2 3 6 7
0
0 0 624 180
6 74LS22
-21 -28 21 -20
3 U3A
-8 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
8745 0 0
2
5.89886e-315 0
0
6 JK RN~
219 702 233 0 6 22
0 9 5 9 7 10 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
9592 0 0
2
5.89886e-315 5.26354e-315
0
6 JK RN~
219 847 235 0 6 22
0 9 3 9 7 11 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
8748 0 0
2
5.89886e-315 0
0
6 JK RN~
219 571 235 0 6 22
0 9 6 9 7 12 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
7168 0 0
2
5.89886e-315 0
0
6 JK RN~
219 426 233 0 6 22
0 9 8 9 7 13 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
631 0 0
2
5.89886e-315 0
0
25
2 2 2 0 0 4224 0 3 8 0 0 3
990 242
990 281
968 281
0 3 3 0 0 4224 0 0 8 14 0 4
775 136
1006 136
1006 293
968 293
0 1 4 0 0 8320 0 0 8 13 0 4
910 128
1025 128
1025 305
968 305
0 1 5 0 0 4224 0 0 3 15 0 3
632 141
990 141
990 206
0 4 6 0 0 4224 0 0 8 16 0 4
486 148
980 148
980 269
968 269
4 0 7 0 0 4096 0 10 0 0 9 2
847 266
847 287
4 0 7 0 0 0 0 9 0 0 9 4
702 264
702 282
703 282
703 287
4 0 7 0 0 0 0 11 0 0 9 2
571 266
571 287
5 4 7 0 0 4224 0 8 12 0 0 3
917 287
426 287
426 264
2 0 6 0 0 0 0 11 0 0 16 3
540 227
480 227
480 216
2 0 3 0 0 0 0 10 0 0 14 3
816 227
767 227
767 216
2 0 5 0 0 0 0 9 0 0 15 3
671 225
631 225
631 218
6 1 4 0 0 0 0 10 4 0 0 5
871 218
910 218
910 128
737 128
737 118
6 1 3 0 0 0 0 9 5 0 0 3
726 216
775 216
775 116
6 1 5 0 0 0 0 11 6 0 0 5
595 218
632 218
632 141
811 141
811 117
6 1 6 0 0 0 0 12 7 0 0 5
450 216
486 216
486 148
845 148
845 116
1 2 8 0 0 4224 0 1 12 0 0 4
255 220
387 220
387 225
395 225
1 0 9 0 0 4096 0 12 0 0 19 2
402 216
363 216
3 0 9 0 0 8192 0 12 0 0 25 3
402 234
363 234
363 155
1 0 9 0 0 0 0 11 0 0 21 2
547 218
523 218
3 0 9 0 0 8192 0 11 0 0 25 3
547 236
523 236
523 155
1 0 9 0 0 0 0 9 0 0 23 2
678 216
661 216
3 0 9 0 0 0 0 9 0 0 25 3
678 234
661 234
661 155
1 0 9 0 0 0 0 10 0 0 25 2
823 218
802 218
3 1 9 0 0 12416 0 10 2 0 0 4
823 236
802 236
802 155
252 155
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
