CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 728 206 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4331 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 745 253 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
787 0 0
2
5.89886e-315 5.26354e-315
0
13 Logic Switch~
5 599 247 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3655 0 0
2
5.89886e-315 5.30499e-315
0
13 Logic Switch~
5 591 203 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6682 0 0
2
5.89886e-315 5.32571e-315
0
13 Logic Switch~
5 468 201 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
582 0 0
2
5.89886e-315 5.34643e-315
0
13 Logic Switch~
5 478 248 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3125 0 0
2
5.89886e-315 5.3568e-315
0
13 Logic Switch~
5 355 207 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5466 0 0
2
5.89886e-315 5.36716e-315
0
13 Logic Switch~
5 354 247 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
52 0 0
2
5.89886e-315 5.37752e-315
0
13 Logic Switch~
5 864 221 0 1 11
0 6
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3898 0 0
2
5.89886e-315 5.38788e-315
0
5 4027~
219 262 243 0 7 32
0 18 15 17 14 19 20 5
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U3B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
9413 0 0
2
5.89886e-315 5.39306e-315
0
5 4027~
219 410 248 0 7 32
0 21 12 16 11 22 17 4
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U3A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
8576 0 0
2
5.89886e-315 5.39824e-315
0
5 4027~
219 531 249 0 7 32
0 23 9 7 10 24 16 3
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
622 0 0
2
5.89886e-315 5.40342e-315
0
5 4027~
219 664 248 0 7 32
0 25 13 6 8 26 7 2
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9152 0 0
2
5.89886e-315 5.4086e-315
0
14 Logic Display~
6 614 105 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
783 0 0
2
5.89886e-315 5.41378e-315
0
14 Logic Display~
6 487 103 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4262 0 0
2
5.89886e-315 5.41896e-315
0
14 Logic Display~
6 372 106 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6121 0 0
2
5.89886e-315 5.42414e-315
0
14 Logic Display~
6 235 105 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3879 0 0
2
5.89886e-315 5.42933e-315
0
16
1 7 2 0 0 4224 0 14 13 0 0 3
614 123
614 212
646 212
1 7 3 0 0 4224 0 15 12 0 0 3
487 121
487 213
513 213
1 7 4 0 0 4224 0 16 11 0 0 3
372 124
372 212
392 212
1 7 5 0 0 4224 0 17 10 0 0 3
235 123
235 207
244 207
1 3 6 0 0 4240 0 9 13 0 0 2
852 221
694 221
6 3 7 0 0 4224 0 13 12 0 0 4
640 230
569 230
569 222
561 222
4 1 8 0 0 4224 0 13 2 0 0 4
694 230
727 230
727 253
733 253
1 2 9 0 0 4224 0 4 12 0 0 4
579 203
567 203
567 213
561 213
4 1 10 0 0 12416 0 12 3 0 0 4
561 231
565 231
565 247
587 247
4 1 11 0 0 8320 0 11 6 0 0 4
440 230
452 230
452 248
466 248
1 2 12 0 0 8320 0 5 11 0 0 4
456 201
448 201
448 212
440 212
1 2 13 0 0 4224 0 1 13 0 0 4
716 206
702 206
702 212
694 212
1 4 14 0 0 4224 0 8 10 0 0 4
342 247
300 247
300 225
292 225
1 2 15 0 0 4224 0 7 10 0 0 2
343 207
292 207
6 3 16 0 0 4224 0 12 11 0 0 6
507 231
456 231
456 224
448 224
448 221
440 221
6 3 17 0 0 4224 0 11 10 0 0 6
386 230
313 230
313 217
300 217
300 216
292 216
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
