CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 169 440 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-42 -9 -35 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 162 259 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-35 -7 -28 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 158 137 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 C
-41 -5 -34 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 156 104 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 D
-38 -4 -31 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1046 408 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1043 265 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1041 104 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1039 45 0 1 2
20 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89774e-315 0
0
9 Inverter~
13 367 331 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
6435 0 0
2
5.89774e-315 0
0
9 Inverter~
13 505 219 0 2 22
0 3 2
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
5283 0 0
2
5.89774e-315 0
0
9 Inverter~
13 333 64 0 2 22
0 13 16
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
6874 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 354 122 0 3 22
0 13 14 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5305 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 661 412 0 3 22
0 3 12 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
34 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 651 326 0 3 22
0 3 11 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
969 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 644 250 0 3 22
0 2 12 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8402 0 0
2
5.89774e-315 0
0
8 2-In OR~
219 351 217 0 3 22
0 13 14 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3751 0 0
2
5.89774e-315 0
0
8 2-In OR~
219 623 132 0 3 22
0 15 2 4
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4292 0 0
2
5.89774e-315 0
0
8 2-In OR~
219 858 431 0 3 22
0 10 9 5
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6118 0 0
2
5.89774e-315 0
0
8 2-In OR~
219 844 283 0 3 22
0 8 7 6
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
34 0 0
2
5.89774e-315 0
0
23
0 2 2 0 0 4096 0 0 17 15 0 3
589 219
589 141
610 141
1 0 3 0 0 4096 0 14 0 0 11 2
627 317
454 317
3 1 4 0 0 4224 0 17 7 0 0 3
656 132
1041 132
1041 122
3 1 5 0 0 4224 0 18 5 0 0 3
891 431
1046 431
1046 426
3 1 6 0 0 4224 0 19 6 0 0 2
877 283
1043 283
3 2 7 0 0 12416 0 14 19 0 0 4
672 326
687 326
687 292
831 292
1 3 8 0 0 4224 0 19 15 0 0 4
831 274
673 274
673 250
665 250
2 1 9 0 0 4224 0 18 1 0 0 2
845 440
181 440
3 1 10 0 0 4224 0 13 18 0 0 4
682 412
837 412
837 422
845 422
2 2 11 0 0 4224 0 14 9 0 0 4
627 335
396 335
396 331
388 331
0 1 3 0 0 4224 0 0 13 16 0 3
454 217
454 403
637 403
0 1 12 0 0 4096 0 0 9 13 0 2
210 331
352 331
0 2 12 0 0 8192 0 0 13 14 0 3
210 259
210 421
637 421
1 2 12 0 0 4224 0 2 15 0 0 2
174 259
620 259
2 1 2 0 0 4224 0 10 15 0 0 4
526 219
612 219
612 241
620 241
3 1 3 0 0 0 0 16 10 0 0 4
384 217
482 217
482 219
490 219
0 1 13 0 0 4096 0 0 16 19 0 3
281 104
281 208
338 208
1 0 13 0 0 4096 0 11 0 0 19 3
318 64
212 64
212 104
1 1 13 0 0 4224 0 4 12 0 0 4
168 104
322 104
322 113
330 113
0 2 14 0 0 8192 0 0 16 22 0 3
190 137
190 226
338 226
1 3 15 0 0 4224 0 17 12 0 0 4
610 123
383 123
383 122
375 122
1 2 14 0 0 4224 0 3 12 0 0 4
170 137
322 137
322 131
330 131
1 2 16 0 0 8320 0 8 11 0 0 5
1039 63
1039 67
362 67
362 64
354 64
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1005 390 1030 414
1013 398 1021 414
1 w
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
996 245 1025 269
1006 253 1014 269
1 x
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
992 99 1021 123
1002 107 1010 123
1 y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
993 39 1022 63
1003 47 1011 63
1 z
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
