CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 214 535 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -14 8 -6
1 A
-34 -6 -27 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42666.9 0
0
13 Logic Switch~
5 216 376 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-36 -5 -29 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
42666.9 0
0
13 Logic Switch~
5 211 259 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-33 -4 -26 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
42666.9 0
0
13 Logic Switch~
5 206 115 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-32 -5 -25 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
42666.9 0
0
14 Logic Display~
6 1129 450 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
42666.9 0
0
14 Logic Display~
6 1123 300 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
42666.9 0
0
14 Logic Display~
6 1113 160 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
42666.9 0
0
14 Logic Display~
6 1108 80 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
42666.9 0
0
8 2-In OR~
219 1040 317 0 3 22
0 17 14 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4747 0 0
2
42666.9 0
0
9 2-In AND~
219 930 273 0 3 22
0 18 4 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
972 0 0
2
42666.9 0
0
8 2-In OR~
219 925 467 0 3 22
0 13 12 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3472 0 0
2
42666.9 0
0
9 2-In AND~
219 761 503 0 3 22
0 10 11 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9998 0 0
2
42666.9 0
0
8 3-In OR~
219 634 495 0 4 22
0 2 3 4 10
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
3536 0 0
2
42666.9 0
0
9 4-In AND~
219 749 431 0 5 22
0 8 6 7 5 13
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U5A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
4597 0 0
2
42666.9 0
0
9 Inverter~
13 729 263 0 2 22
0 9 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3835 0 0
2
42666.9 0
0
9 2-In AND~
219 741 354 0 3 22
0 9 6 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3670 0 0
2
42666.9 0
0
8 2-In OR~
219 585 261 0 3 22
0 3 2 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5616 0 0
2
42666.9 0
0
6 74136~
219 593 188 0 3 22
0 2 3 19
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
42666.9 0
0
9 Inverter~
13 421 535 0 2 22
0 5 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
317 0 0
2
42666.9 0
0
9 Inverter~
13 408 376 0 2 22
0 4 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3108 0 0
2
42666.9 0
0
9 Inverter~
13 400 259 0 2 22
0 3 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4299 0 0
2
42666.9 0
0
9 Inverter~
13 396 151 0 2 22
0 2 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9672 0 0
2
42666.9 0
0
30
0 1 2 0 0 4096 0 0 13 29 0 3
357 151
357 486
621 486
0 2 3 0 0 8320 0 0 13 26 0 3
334 259
334 495
622 495
0 3 4 0 0 8192 0 0 13 25 0 3
321 376
321 504
621 504
4 0 5 0 0 4224 0 14 0 0 24 3
725 445
312 445
312 535
0 2 6 0 0 8192 0 0 14 8 0 3
631 376
631 427
725 427
2 3 7 0 0 8320 0 21 14 0 0 4
421 259
568 259
568 436
725 436
2 1 8 0 0 4224 0 22 14 0 0 4
417 151
699 151
699 418
725 418
2 2 6 0 0 4224 0 20 16 0 0 4
429 376
709 376
709 363
717 363
2 0 4 0 0 4224 0 10 0 0 25 3
906 282
280 282
280 376
0 1 9 0 0 4096 0 0 16 20 0 3
659 261
659 345
717 345
4 1 10 0 0 4224 0 13 12 0 0 4
667 495
729 495
729 494
737 494
2 2 11 0 0 4224 0 19 12 0 0 4
442 535
729 535
729 512
737 512
3 2 12 0 0 4224 0 12 11 0 0 4
782 503
904 503
904 476
912 476
5 1 13 0 0 4224 0 14 11 0 0 4
770 431
904 431
904 458
912 458
3 2 14 0 0 4224 0 16 9 0 0 4
762 354
1019 354
1019 326
1027 326
3 1 15 0 0 4224 0 11 5 0 0 3
958 467
1129 467
1129 468
3 1 16 0 0 4224 0 9 6 0 0 3
1073 317
1123 317
1123 318
3 1 17 0 0 4224 0 10 9 0 0 4
951 273
1019 273
1019 308
1027 308
2 1 18 0 0 4224 0 15 10 0 0 4
750 263
898 263
898 264
906 264
3 1 9 0 0 4224 0 17 15 0 0 4
618 261
706 261
706 263
714 263
0 2 2 0 0 0 0 0 17 30 0 3
455 115
455 270
572 270
1 0 3 0 0 0 0 17 0 0 23 3
572 252
525 252
525 197
2 0 3 0 0 0 0 18 0 0 26 3
577 197
293 197
293 259
1 1 5 0 0 0 0 1 19 0 0 2
226 535
406 535
1 1 4 0 0 0 0 2 20 0 0 2
228 376
393 376
1 1 3 0 0 0 0 3 21 0 0 2
223 259
385 259
3 1 19 0 0 4224 0 18 7 0 0 3
626 188
1113 188
1113 178
1 0 2 0 0 0 0 18 0 0 30 3
577 179
545 179
545 115
1 0 2 0 0 0 0 22 0 0 30 3
381 151
280 151
280 115
1 1 2 0 0 4224 0 4 8 0 0 3
218 115
1108 115
1108 98
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1083 442 1120 466
1093 450 1109 466
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1083 289 1120 313
1093 297 1109 313
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1067 159 1104 183
1077 167 1093 183
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1064 88 1101 112
1074 96 1090 112
2 S4
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
