CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
44
13 Logic Switch~
5 497 606 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 181 315 0 1 11
0 39
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 365 190 0 1 11
0 42
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 E
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 363 131 0 1 11
0 43
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 361 64 0 1 11
0 44
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 182 262 0 1 11
0 40
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 176 204 0 1 11
0 41
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89886e-315 0
0
7 74LS138
19 672 138 0 14 29
0 44 43 42 38 2 2 27 28 29
30 31 32 33 34
0
0 0 5088 0
6 74F138
-21 -61 21 -53
2 U2
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7361 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 999 519 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L24
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89886e-315 5.37752e-315
0
14 Logic Display~
6 967 519 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L25
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89886e-315 5.36716e-315
0
14 Logic Display~
6 936 521 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L26
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89886e-315 5.3568e-315
0
14 Logic Display~
6 908 520 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L27
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89886e-315 5.34643e-315
0
14 Logic Display~
6 879 519 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L28
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 849 518 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L29
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 816 519 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L30
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 791 520 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L31
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 995 369 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89886e-315 5.37752e-315
0
14 Logic Display~
6 968 369 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89886e-315 5.36716e-315
0
14 Logic Display~
6 938 369 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89886e-315 5.3568e-315
0
14 Logic Display~
6 909 369 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89886e-315 5.34643e-315
0
14 Logic Display~
6 878 369 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 848 370 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 818 371 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L22
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 790 372 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L23
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 1018 218 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89886e-315 5.37752e-315
0
14 Logic Display~
6 981 218 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89886e-315 5.36716e-315
0
14 Logic Display~
6 944 219 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89886e-315 5.3568e-315
0
14 Logic Display~
6 909 218 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89886e-315 5.34643e-315
0
14 Logic Display~
6 875 220 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 846 219 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 817 218 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 782 218 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 845 64 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89886e-315 5.37752e-315
0
14 Logic Display~
6 821 63 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89886e-315 5.36716e-315
0
14 Logic Display~
6 782 63 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.89886e-315 5.3568e-315
0
14 Logic Display~
6 1030 65 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.89886e-315 5.34643e-315
0
14 Logic Display~
6 885 65 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 921 64 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 960 65 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 999 66 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89886e-315 0
0
7 74LS138
19 674 572 0 14 29
0 44 43 42 35 2 2 3 4 5
6 7 8 9 10
0
0 0 5088 0
6 74F138
-21 -61 21 -53
2 U5
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
5.89886e-315 0
0
7 74LS138
19 674 443 0 14 29
0 44 43 42 36 2 2 11 12 13
14 15 16 17 18
0
0 0 5088 0
6 74F138
-21 -61 21 -53
2 U4
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3171 0 0
2
5.89886e-315 0
0
7 74LS138
19 673 290 0 14 29
0 44 43 42 37 2 2 19 20 21
22 23 24 25 26
0
0 0 5088 0
6 74F138
-21 -61 21 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4139 0 0
2
5.89886e-315 0
0
4 4555
219 300 253 0 7 32
0 41 40 39 38 37 36 35
0
0 0 4832 0
4 4555
-14 -60 14 -52
3 U1A
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 3 2 1 4 5 6 7 3 2
1 4 5 6 7 13 14 15 12 11
10 9 0 0 0 0 0 0 0 0
0 19 0
65 0 0 0 2 1 1 0
1 U
6435 0 0
2
5.89886e-315 0
0
59
6 0 2 0 0 4096 0 41 0 0 8 2
636 608
629 608
5 0 2 0 0 0 0 41 0 0 8 2
636 599
629 599
6 0 2 0 0 0 0 42 0 0 8 2
636 479
629 479
5 0 2 0 0 0 0 42 0 0 8 2
636 470
629 470
6 0 2 0 0 0 0 43 0 0 8 2
635 326
629 326
5 0 2 0 0 0 0 43 0 0 8 2
635 317
629 317
6 0 2 0 0 0 0 8 0 0 8 2
634 174
629 174
1 5 2 0 0 8320 0 1 8 0 0 6
509 606
629 606
629 608
629 608
629 165
634 165
7 1 3 0 0 4224 0 41 16 0 0 3
712 545
791 545
791 538
8 1 4 0 0 4224 0 41 15 0 0 3
712 554
816 554
816 537
9 1 5 0 0 4224 0 41 14 0 0 3
712 563
849 563
849 536
1 10 6 0 0 8320 0 13 41 0 0 3
879 537
879 572
712 572
11 1 7 0 0 4224 0 41 12 0 0 3
712 581
908 581
908 538
12 1 8 0 0 4224 0 41 11 0 0 3
712 590
936 590
936 539
13 1 9 0 0 4224 0 41 10 0 0 3
712 599
967 599
967 537
14 1 10 0 0 4224 0 41 9 0 0 3
712 608
999 608
999 537
7 1 11 0 0 4224 0 42 24 0 0 3
712 416
790 416
790 390
8 1 12 0 0 4224 0 42 23 0 0 3
712 425
818 425
818 389
9 1 13 0 0 4224 0 42 22 0 0 3
712 434
848 434
848 388
10 1 14 0 0 4224 0 42 21 0 0 3
712 443
878 443
878 387
11 1 15 0 0 4224 0 42 20 0 0 3
712 452
909 452
909 387
12 1 16 0 0 4224 0 42 19 0 0 3
712 461
938 461
938 387
13 1 17 0 0 4224 0 42 18 0 0 3
712 470
968 470
968 387
14 1 18 0 0 4224 0 42 17 0 0 3
712 479
995 479
995 387
1 7 19 0 0 8320 0 32 43 0 0 3
782 236
782 263
711 263
8 1 20 0 0 4224 0 43 31 0 0 3
711 272
817 272
817 236
9 1 21 0 0 4224 0 43 30 0 0 3
711 281
846 281
846 237
10 1 22 0 0 4224 0 43 29 0 0 3
711 290
875 290
875 238
11 1 23 0 0 4224 0 43 28 0 0 3
711 299
909 299
909 236
12 1 24 0 0 4224 0 43 27 0 0 3
711 308
944 308
944 237
13 1 25 0 0 4224 0 43 26 0 0 3
711 317
981 317
981 236
14 1 26 0 0 4224 0 43 25 0 0 3
711 326
1018 326
1018 236
7 1 27 0 0 4224 0 8 35 0 0 3
710 111
782 111
782 81
8 1 28 0 0 4224 0 8 34 0 0 3
710 120
821 120
821 81
9 1 29 0 0 4224 0 8 33 0 0 3
710 129
845 129
845 82
10 1 30 0 0 4224 0 8 37 0 0 3
710 138
885 138
885 83
11 1 31 0 0 4224 0 8 38 0 0 3
710 147
921 147
921 82
12 1 32 0 0 4224 0 8 39 0 0 3
710 156
960 156
960 83
13 1 33 0 0 4224 0 8 40 0 0 3
710 165
999 165
999 84
14 1 34 0 0 4240 0 8 36 0 0 3
710 174
1030 174
1030 83
7 4 35 0 0 12416 0 44 41 0 0 5
332 226
332 211
597 211
597 590
642 590
6 4 36 0 0 4224 0 44 42 0 0 4
332 235
608 235
608 461
642 461
5 4 37 0 0 4224 0 44 43 0 0 4
332 244
615 244
615 308
641 308
4 4 38 0 0 4224 0 44 8 0 0 4
332 253
621 253
621 156
640 156
1 3 39 0 0 4224 0 2 44 0 0 3
193 315
262 315
262 253
1 2 40 0 0 4224 0 6 44 0 0 4
194 262
253 262
253 235
268 235
1 1 41 0 0 4224 0 7 44 0 0 4
188 204
254 204
254 226
268 226
0 3 42 0 0 4096 0 0 41 49 0 3
585 433
585 563
642 563
0 3 42 0 0 4096 0 0 42 50 0 3
585 281
585 434
642 434
0 3 42 0 0 0 0 0 43 51 0 3
585 129
585 281
641 281
1 3 42 0 0 4224 0 3 8 0 0 4
377 190
585 190
585 129
640 129
0 2 43 0 0 4096 0 0 41 53 0 3
563 425
563 554
642 554
0 2 43 0 0 4096 0 0 42 54 0 3
563 271
563 425
642 425
0 2 43 0 0 0 0 0 43 55 0 3
563 120
563 272
641 272
1 2 43 0 0 4224 0 4 8 0 0 4
375 131
563 131
563 120
640 120
0 1 44 0 0 4096 0 0 41 57 0 3
525 416
525 545
642 545
0 1 44 0 0 4224 0 0 42 58 0 3
525 263
525 416
642 416
0 1 44 0 0 0 0 0 43 59 0 3
525 110
525 263
641 263
1 1 44 0 0 0 0 5 8 0 0 4
373 64
525 64
525 111
640 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
