CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
19
14 Logic Display~
6 773 238 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5130 0 0
2
43556.7 0
0
14 Logic Display~
6 765 76 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
43556.7 0
0
14 Logic Display~
6 777 340 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3124 0 0
2
43556.7 0
0
13 Logic Switch~
5 243 441 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 G1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3421 0 0
2
43556.7 0
0
13 Logic Switch~
5 246 406 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 P1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8157 0 0
2
43556.7 0
0
13 Logic Switch~
5 242 322 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 P2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
43556.7 0
0
13 Logic Switch~
5 242 481 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 C1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
43556.7 0
0
13 Logic Switch~
5 240 357 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 G2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
43556.7 0
0
13 Logic Switch~
5 240 197 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 P3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
43556.7 0
0
13 Logic Switch~
5 242 236 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 G3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43556.7 0
0
8 2-In OR~
219 574 406 0 1 22
0 0
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3472 0 0
2
43556.7 0
0
8 3-In OR~
219 573 285 0 1 22
0 0
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
9998 0 0
2
43556.7 0
0
8 4-In OR~
219 577 131 0 1 22
0 0
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
3536 0 0
2
43556.7 0
0
9 2-In AND~
219 406 397 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4597 0 0
2
43556.7 0
0
5 7415~
219 403 268 0 1 22
0 0
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
3835 0 0
2
43556.7 0
0
5 7415~
219 398 138 0 1 22
0 0
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
3670 0 0
2
43556.7 0
0
9 4-In AND~
219 397 85 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
5616 0 0
2
43556.7 0
0
9 2-In AND~
219 400 188 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
43556.7 0
0
9 2-In AND~
219 404 313 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
317 0 0
2
43556.7 0
0
28
1 0 0 0 0 0 0 14 0 0 13 2
382 388
361 388
1 0 0 0 0 0 0 19 0 0 9 2
380 304
347 304
3 0 0 0 0 0 0 15 0 0 11 2
379 277
305 277
2 0 0 0 0 0 0 15 0 0 10 2
379 268
275 268
1 0 0 0 0 0 0 15 0 0 13 2
379 259
361 259
0 1 0 0 0 0 0 0 18 16 0 3
323 357
323 179
376 179
3 0 0 0 0 0 0 16 0 0 12 2
374 147
337 147
2 0 0 0 0 0 0 16 0 0 11 2
374 138
305 138
0 1 0 0 0 0 0 0 16 15 0 3
347 441
347 129
374 129
0 1 0 0 0 0 0 0 17 14 0 3
275 406
275 72
373 72
0 2 0 0 0 0 0 0 17 17 0 3
305 322
305 81
373 81
0 3 0 0 0 0 0 0 17 19 0 3
337 197
337 90
373 90
1 4 0 0 0 0 0 7 17 0 0 4
254 481
361 481
361 99
373 99
1 2 0 0 0 0 0 5 14 0 0 2
258 406
382 406
1 2 0 0 0 0 0 4 11 0 0 4
255 441
542 441
542 415
561 415
1 3 0 0 0 0 0 8 12 0 0 4
252 357
542 357
542 294
560 294
1 2 0 0 0 0 0 6 19 0 0 2
254 322
380 322
1 4 0 0 0 0 0 10 13 0 0 4
254 236
541 236
541 145
560 145
1 2 0 0 0 0 0 9 18 0 0 2
252 197
376 197
3 1 0 0 0 0 0 14 11 0 0 2
427 397
561 397
3 2 0 0 0 0 0 19 12 0 0 4
425 313
524 313
524 285
561 285
4 1 0 0 0 0 0 15 12 0 0 4
424 268
524 268
524 276
560 276
3 3 0 0 0 0 0 18 13 0 0 4
421 188
530 188
530 136
560 136
4 2 0 0 0 0 0 16 13 0 0 4
419 138
523 138
523 127
560 127
5 1 0 0 0 0 0 17 13 0 0 4
418 85
523 85
523 118
560 118
1 3 0 0 0 0 0 3 11 0 0 3
777 358
777 406
607 406
1 4 0 0 0 0 0 1 12 0 0 3
773 256
773 285
606 285
5 1 0 0 0 0 0 13 2 0 0 3
610 131
765 131
765 94
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
