CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 833 306 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-6 -14 8 -6
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5789 0 0
2
5.89864e-315 0
0
13 Logic Switch~
5 968 254 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7328 0 0
2
5.89864e-315 0
0
14 Logic Display~
6 804 74 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4799 0 0
2
5.89864e-315 0
0
14 Logic Display~
6 636 75 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9196 0 0
2
5.89864e-315 0
0
14 Logic Display~
6 511 71 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3857 0 0
2
5.89864e-315 0
0
14 Logic Display~
6 399 74 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7125 0 0
2
5.89864e-315 0
0
5 4049~
219 850 254 0 2 22
0 2 7
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U4A
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
3641 0 0
2
5.89864e-315 0
0
9 2-In AND~
219 323 269 0 3 22
0 3 8 12
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 3 0
1 U
9821 0 0
2
5.89864e-315 0
0
9 2-In AND~
219 433 281 0 3 22
0 4 9 8
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3187 0 0
2
5.89864e-315 0
0
9 2-In AND~
219 560 289 0 3 22
0 5 10 9
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
762 0 0
2
5.89864e-315 0
0
9 2-In AND~
219 702 297 0 3 22
0 6 11 10
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
39 0 0
2
5.89864e-315 0
0
5 4027~
219 386 227 0 7 32
0 13 8 7 8 14 15 3
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U2B
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9450 0 0
2
5.89864e-315 0
0
5 4027~
219 500 230 0 7 32
0 16 9 7 9 17 18 4
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U2A
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3236 0 0
2
5.89864e-315 0
0
5 4027~
219 623 228 0 7 32
0 19 10 7 10 20 21 5
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U1B
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3321 0 0
2
5.89864e-315 0
0
5 4027~
219 791 230 0 7 32
0 22 11 7 11 23 24 6
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U1A
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
8879 0 0
2
5.89864e-315 0
0
25
1 1 2 0 0 4224 0 7 2 0 0 2
871 254
956 254
1 0 3 0 0 4096 0 6 0 0 10 2
399 92
399 172
1 0 4 0 0 4096 0 5 0 0 14 3
511 89
511 173
513 173
1 0 5 0 0 4096 0 4 0 0 18 2
636 93
636 171
1 0 6 0 0 4096 0 3 0 0 22 2
804 92
804 173
3 0 7 0 0 4096 0 13 0 0 9 4
504 231
504 249
505 249
505 254
3 0 7 0 0 4096 0 14 0 0 9 2
627 229
627 254
3 0 7 0 0 0 0 15 0 0 9 4
795 231
795 249
796 249
796 254
3 2 7 0 0 8320 0 12 7 0 0 3
390 228
390 254
835 254
7 1 3 0 0 12416 0 12 8 0 0 5
399 180
399 170
352 170
352 260
343 260
4 0 8 0 0 4096 0 12 0 0 13 2
381 228
381 281
2 0 8 0 0 0 0 12 0 0 13 2
399 228
399 281
3 2 8 0 0 4224 0 9 8 0 0 4
408 281
352 281
352 278
343 278
7 1 4 0 0 12416 0 13 9 0 0 5
513 183
513 173
462 173
462 272
453 272
4 0 9 0 0 4096 0 13 0 0 17 2
495 231
495 289
2 0 9 0 0 0 0 13 0 0 17 2
513 231
513 289
3 2 9 0 0 4224 0 10 9 0 0 4
535 289
462 289
462 290
453 290
7 1 5 0 0 12416 0 14 10 0 0 5
636 181
636 171
589 171
589 280
580 280
4 0 10 0 0 4096 0 14 0 0 21 2
618 229
618 297
2 0 10 0 0 0 0 14 0 0 21 2
636 229
636 297
3 2 10 0 0 4224 0 11 10 0 0 4
677 297
589 297
589 298
580 298
7 1 6 0 0 12416 0 15 11 0 0 5
804 183
804 173
731 173
731 288
722 288
4 0 11 0 0 4096 0 15 0 0 25 2
786 231
786 306
2 0 11 0 0 0 0 15 0 0 25 2
804 231
804 306
2 1 11 0 0 4224 0 11 1 0 0 2
722 306
821 306
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
