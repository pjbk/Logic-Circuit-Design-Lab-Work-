CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 361 309 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-56 -10 -49 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7311 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 355 184 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-51 -5 -44 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3409 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 810 258 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3526 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 806 164 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4129 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 631 280 0 3 22
0 5 4 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6278 0 0
2
5.89774e-315 0
0
6 74136~
219 565 187 0 3 22
0 5 4 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3482 0 0
2
5.89774e-315 0
0
6
3 1 2 0 0 4224 0 5 3 0 0 3
652 280
810 280
810 276
3 1 3 0 0 4224 0 6 4 0 0 3
598 187
806 187
806 182
2 0 4 0 0 4096 0 5 0 0 5 2
607 289
541 289
1 0 5 0 0 4224 0 5 0 0 6 3
607 271
418 271
418 184
1 2 4 0 0 4224 0 1 6 0 0 4
373 309
541 309
541 196
549 196
1 1 5 0 0 0 0 2 6 0 0 4
367 184
541 184
541 178
549 178
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
715 243 776 265
725 250 765 266
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
717 160 760 182
726 167 750 183
3 sum
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
