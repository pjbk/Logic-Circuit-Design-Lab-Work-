CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 108 144 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 x
-42 -6 -35 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
43549.9 2
0
13 Logic Switch~
5 106 249 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 y
-39 -12 -32 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3674 0 0
2
43549.9 1
0
13 Logic Switch~
5 100 419 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 bin
-48 -9 -27 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5697 0 0
2
43549.9 0
0
9 Inverter~
13 727 167 0 2 22
0 4 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3805 0 0
2
43549.9 0
0
9 Inverter~
13 138 144 0 2 22
0 13 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
5219 0 0
2
43549.9 0
0
6 74136~
219 648 167 0 3 22
0 10 8 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3795 0 0
2
43549.9 11
0
6 74136~
219 297 154 0 3 22
0 3 12 10
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3637 0 0
2
43549.9 10
0
9 2-In AND~
219 323 333 0 3 22
0 12 11 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3226 0 0
2
43549.9 9
0
9 2-In AND~
219 764 257 0 3 22
0 9 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6966 0 0
2
43549.9 8
0
8 2-In OR~
219 849 312 0 3 22
0 6 7 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9796 0 0
2
43549.9 7
0
14 Logic Display~
6 1075 149 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
43549.9 6
0
14 Logic Display~
6 1063 294 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
43549.9 5
0
9 Inverter~
13 200 342 0 2 22
0 3 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3716 0 0
2
43549.9 4
0
9 Inverter~
13 667 248 0 2 22
0 10 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4797 0 0
2
43549.9 3
0
16
2 1 2 0 0 4240 0 4 11 0 0 2
748 167
1075 167
2 1 3 0 0 4112 0 5 7 0 0 4
159 144
273 144
273 145
281 145
3 1 4 0 0 4240 0 6 4 0 0 2
681 167
712 167
3 1 5 0 0 4240 0 10 12 0 0 2
882 312
1063 312
3 1 6 0 0 8336 0 9 10 0 0 4
785 257
828 257
828 303
836 303
3 2 7 0 0 4240 0 8 10 0 0 4
344 333
821 333
821 321
836 321
2 0 8 0 0 4112 0 9 0 0 10 2
740 266
624 266
2 1 9 0 0 4240 0 14 9 0 0 2
688 248
740 248
0 1 10 0 0 8208 0 0 14 11 0 3
431 154
431 248
652 248
1 2 8 0 0 4240 0 3 6 0 0 4
112 419
624 419
624 176
632 176
3 1 10 0 0 4240 0 7 6 0 0 4
330 154
624 154
624 158
632 158
0 1 3 0 0 4240 0 0 13 2 0 3
165 144
165 342
185 342
2 2 11 0 0 4240 0 13 8 0 0 2
221 342
299 342
1 0 12 0 0 8208 0 8 0 0 15 4
299 324
288 324
288 249
273 249
1 2 12 0 0 4240 0 2 7 0 0 4
118 249
273 249
273 163
281 163
1 1 13 0 0 4240 0 1 5 0 0 2
120 144
123 144
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1025 139 1054 163
1035 147 1043 163
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1004 278 1057 302
1014 286 1046 302
4 bout
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
