CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 80 152 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44175.5 0
0
13 Logic Switch~
5 81 223 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
44175.5 1
0
9 Inverter~
13 593 446 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4597 0 0
2
44175.5 2
0
9 Inverter~
13 470 303 0 2 22
0 6 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3835 0 0
2
44175.5 3
0
14 Logic Display~
6 649 106 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
44175.5 4
0
14 Logic Display~
6 696 106 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44175.5 5
0
14 Logic Display~
6 737 105 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
44175.5 6
0
5 7415~
219 499 416 0 4 22
0 7 5 4 3
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
317 0 0
2
44175.5 7
0
6 JK RN~
219 601 231 0 6 22
0 9 6 9 2 10 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
3108 0 0
2
44175.5 8
0
6 JK RN~
219 404 229 0 6 22
0 9 4 9 2 11 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
4299 0 0
2
44175.5 9
0
6 JK RN~
219 229 230 0 6 22
0 9 8 9 2 12 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9672 0 0
2
44175.5 10
0
20
0 4 2 0 0 4096 0 0 10 2 0 2
404 287
404 260
0 4 2 0 0 4224 0 0 11 3 0 3
618 287
229 287
229 261
2 4 2 0 0 0 0 3 9 0 0 5
614 446
618 446
618 270
601 270
601 262
4 1 3 0 0 4224 0 8 3 0 0 4
520 416
570 416
570 446
578 446
0 3 4 0 0 4224 0 0 8 13 0 3
263 213
263 425
475 425
2 2 5 0 0 8320 0 4 8 0 0 6
491 303
495 303
495 392
470 392
470 416
475 416
0 1 6 0 0 4096 0 0 4 12 0 3
441 212
441 303
455 303
0 1 7 0 0 8320 0 0 8 11 0 5
664 214
664 396
467 396
467 407
475 407
0 1 4 0 0 8336 0 0 7 13 0 4
301 213
301 182
737 182
737 123
0 1 6 0 0 8320 0 0 6 12 0 4
499 212
499 197
696 197
696 124
6 1 7 0 0 0 0 9 5 0 0 5
625 214
664 214
664 214
649 214
649 124
6 2 6 0 0 128 0 10 9 0 0 4
428 212
557 212
557 223
570 223
6 2 4 0 0 0 0 11 10 0 0 4
253 213
365 213
365 221
373 221
1 2 8 0 0 4224 0 2 11 0 0 4
93 223
190 223
190 222
198 222
3 0 9 0 0 8192 0 11 0 0 20 3
205 231
169 231
169 152
1 0 9 0 0 0 0 11 0 0 20 3
205 213
193 213
193 152
3 0 9 0 0 0 0 10 0 0 20 3
380 230
346 230
346 152
1 0 9 0 0 0 0 10 0 0 20 3
380 212
369 212
369 152
3 0 9 0 0 8192 0 9 0 0 20 3
577 232
541 232
541 152
1 1 9 0 0 4224 0 1 9 0 0 4
92 152
562 152
562 214
577 214
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
