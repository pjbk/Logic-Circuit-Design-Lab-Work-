CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 354 424 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3723 0 0
2
43809.8 0
0
13 Logic Switch~
5 350 330 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3440 0 0
2
43809.8 0
0
13 Logic Switch~
5 348 270 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6263 0 0
2
43809.8 0
0
13 Logic Switch~
5 346 225 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4900 0 0
2
43809.8 0
0
13 Logic Switch~
5 336 161 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8783 0 0
2
43809.8 0
0
13 Logic Switch~
5 336 122 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3221 0 0
2
43809.8 0
0
14 Logic Display~
6 639 356 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3215 0 0
2
43809.8 0
0
9 2-In NOR~
219 553 378 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7903 0 0
2
43809.8 0
0
9 2-In NOR~
219 465 415 0 3 22
0 2 2 5
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7121 0 0
2
43809.8 0
0
9 2-In NOR~
219 464 339 0 3 22
0 3 3 6
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4484 0 0
2
43809.8 0
0
14 Logic Display~
6 630 229 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5996 0 0
2
43809.8 0
0
10 2-In NAND~
219 554 247 0 3 22
0 8 8 7
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7804 0 0
2
43809.8 0
0
10 2-In NAND~
219 469 245 0 3 22
0 10 9 8
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5523 0 0
2
43809.8 0
0
14 Logic Display~
6 621 116 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3330 0 0
2
43809.8 0
0
9 2-In AND~
219 490 139 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3465 0 0
2
43809.8 0
0
15
0 1 2 0 0 8192 0 0 9 4 0 3
420 424
420 406
452 406
0 2 3 0 0 8192 0 0 10 3 0 3
418 330
418 348
451 348
1 1 3 0 0 4224 0 2 10 0 0 2
362 330
451 330
1 2 2 0 0 4224 0 1 9 0 0 2
366 424
452 424
3 1 4 0 0 4240 0 8 7 0 0 3
592 378
639 378
639 374
3 2 5 0 0 4224 0 9 8 0 0 4
504 415
532 415
532 387
540 387
3 1 6 0 0 8320 0 10 8 0 0 4
503 339
532 339
532 369
540 369
3 1 7 0 0 4224 0 12 11 0 0 2
581 247
630 247
0 2 8 0 0 4096 0 0 12 10 0 3
519 240
519 256
530 256
3 1 8 0 0 4224 0 13 12 0 0 6
496 245
519 245
519 240
521 240
521 238
530 238
1 2 9 0 0 4224 0 3 13 0 0 4
360 270
437 270
437 254
445 254
1 1 10 0 0 4224 0 4 13 0 0 4
358 225
437 225
437 236
445 236
3 1 11 0 0 4224 0 15 14 0 0 3
511 139
621 139
621 134
1 2 12 0 0 4224 0 5 15 0 0 4
348 161
432 161
432 148
466 148
1 1 13 0 0 4224 0 6 15 0 0 4
348 122
432 122
432 130
466 130
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
99 352 336 376
109 360 325 376
27 AND gate with Universal NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
90 232 335 256
100 240 324 256
28 AND gate with Universal NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
130 125 263 149
140 133 252 149
14 Basic AND gate
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
