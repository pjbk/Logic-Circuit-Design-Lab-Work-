CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 342 201 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89766e-315 0
0
13 Logic Switch~
5 371 164 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89766e-315 0
0
14 Logic Display~
6 665 312 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.89766e-315 0
0
14 Logic Display~
6 664 205 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.89766e-315 0
0
14 Logic Display~
6 665 148 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89766e-315 0
0
10 2-In NAND~
219 564 334 0 3 22
0 6 7 2
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5572 0 0
2
5.89766e-315 0
0
10 2-In NAND~
219 437 375 0 3 22
0 9 10 7
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
5.89766e-315 0
0
10 2-In NAND~
219 438 303 0 3 22
0 8 8 6
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
5.89766e-315 0
0
9 2-In NOR~
219 556 225 0 3 22
0 5 5 3
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
5.89766e-315 0
0
9 2-In NOR~
219 430 225 0 3 22
0 8 9 5
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.89766e-315 0
0
8 2-In OR~
219 431 174 0 3 22
0 8 9 4
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
5.89766e-315 0
0
15
3 1 2 0 0 4224 0 6 3 0 0 3
591 334
665 334
665 330
3 1 3 0 0 4240 0 9 4 0 0 3
595 225
664 225
664 223
3 1 4 0 0 4224 0 11 5 0 0 3
464 174
665 174
665 166
0 2 5 0 0 8192 0 0 9 5 0 3
522 225
522 234
543 234
3 1 5 0 0 4224 0 10 9 0 0 4
469 225
535 225
535 216
543 216
3 1 6 0 0 4224 0 8 6 0 0 4
465 303
532 303
532 325
540 325
3 2 7 0 0 4224 0 7 6 0 0 4
464 375
532 375
532 343
540 343
1 2 8 0 0 8192 0 8 8 0 0 4
414 294
406 294
406 312
414 312
0 1 9 0 0 8320 0 0 7 12 0 4
380 234
400 234
400 366
413 366
0 2 10 0 0 4224 0 0 7 0 0 3
405 366
405 384
413 384
0 1 8 0 0 4224 0 0 8 13 0 3
410 216
410 294
414 294
0 2 9 0 0 0 0 0 10 14 0 3
380 201
380 234
417 234
1 1 8 0 0 0 0 2 10 0 0 4
383 164
404 164
404 216
417 216
1 2 9 0 0 0 0 1 11 0 0 4
354 201
410 201
410 183
418 183
1 1 8 0 0 0 0 2 11 0 0 4
383 164
410 164
410 165
418 165
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
