CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 312 242 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 379 145 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
5.89886e-315 5.26354e-315
0
13 Logic Switch~
5 381 181 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3751 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 379 117 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4292 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 378 77 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6118 0 0
2
5.89886e-315 0
0
9 Inverter~
13 423 181 0 2 22
0 3 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
34 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 926 74 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
5.89886e-315 5.37752e-315
0
14 Logic Display~
6 948 76 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
5.89886e-315 5.36716e-315
0
14 Logic Display~
6 971 75 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
5.89886e-315 5.3568e-315
0
14 Logic Display~
6 993 77 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
5.89886e-315 5.34643e-315
0
14 Logic Display~
6 1083 77 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 1038 76 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 1016 74 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 1061 75 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 800 78 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
5.89886e-315 5.32571e-315
0
14 Logic Display~
6 822 80 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
5.89886e-315 5.30499e-315
0
14 Logic Display~
6 867 81 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.89886e-315 5.26354e-315
0
14 Logic Display~
6 845 79 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 777 81 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 755 79 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 732 80 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 710 78 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.89886e-315 0
0
7 74LS138
19 605 299 0 14 29
0 21 22 23 3 2 2 12 11 10
9 8 7 6 5
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
5.89886e-315 0
0
7 74LS138
19 604 156 0 14 29
0 21 22 23 4 2 2 20 19 18
17 16 15 14 13
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
631 0 0
2
5.89886e-315 0
0
29
6 0 2 0 0 4096 0 23 0 0 2 3
567 335
430 335
430 326
5 0 2 0 0 4224 0 23 0 0 4 3
567 326
418 326
418 242
6 0 2 0 0 0 0 24 0 0 4 2
566 192
448 192
5 1 2 0 0 0 0 24 1 0 0 4
566 183
448 183
448 242
324 242
4 0 3 0 0 4224 0 23 0 0 6 3
573 317
399 317
399 181
1 1 3 0 0 0 0 3 6 0 0 2
393 181
408 181
2 4 4 0 0 4224 0 6 24 0 0 4
444 181
558 181
558 174
572 174
1 14 5 0 0 8320 0 11 23 0 0 3
1083 95
1083 335
643 335
13 1 6 0 0 4224 0 23 14 0 0 3
643 326
1061 326
1061 93
1 12 7 0 0 8320 0 12 23 0 0 3
1038 94
1038 317
643 317
1 11 8 0 0 8320 0 13 23 0 0 3
1016 92
1016 308
643 308
10 1 9 0 0 4224 0 23 10 0 0 3
643 299
993 299
993 95
9 1 10 0 0 4224 0 23 9 0 0 3
643 290
971 290
971 93
8 1 11 0 0 4224 0 23 8 0 0 3
643 281
948 281
948 94
7 1 12 0 0 4224 0 23 7 0 0 3
643 272
926 272
926 92
14 1 13 0 0 4224 0 24 17 0 0 3
642 192
867 192
867 99
13 1 14 0 0 4224 0 24 18 0 0 3
642 183
845 183
845 97
12 1 15 0 0 4224 0 24 16 0 0 3
642 174
822 174
822 98
11 1 16 0 0 4224 0 24 15 0 0 3
642 165
800 165
800 96
10 1 17 0 0 4224 0 24 19 0 0 3
642 156
777 156
777 99
9 1 18 0 0 4224 0 24 20 0 0 3
642 147
755 147
755 97
8 1 19 0 0 4224 0 24 21 0 0 3
642 138
732 138
732 98
7 1 20 0 0 4224 0 24 22 0 0 3
642 129
710 129
710 96
1 0 21 0 0 8320 0 23 0 0 27 3
573 272
514 272
514 77
2 0 22 0 0 8192 0 23 0 0 28 3
573 281
483 281
483 117
3 0 23 0 0 8192 0 23 0 0 29 3
573 290
452 290
452 145
1 1 21 0 0 0 0 5 24 0 0 4
390 77
553 77
553 129
572 129
1 2 22 0 0 4224 0 4 24 0 0 4
391 117
558 117
558 138
572 138
1 3 23 0 0 4224 0 2 24 0 0 4
391 145
558 145
558 147
572 147
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
277 246 362 270
287 254 351 270
8 Always 0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
