CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 288 479 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
44173.5 0
0
13 Logic Switch~
5 287 436 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 D6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
44173.5 0
0
13 Logic Switch~
5 286 397 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
44173.5 0
0
13 Logic Switch~
5 286 359 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9442 0 0
2
44173.5 0
0
13 Logic Switch~
5 287 322 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9424 0 0
2
44173.5 0
0
13 Logic Switch~
5 286 285 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 D2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9968 0 0
2
44173.5 0
0
13 Logic Switch~
5 285 243 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9281 0 0
2
44173.5 0
0
13 Logic Switch~
5 286 200 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -17 8 -9
2 D0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -1 0
1 V
8464 0 0
2
44173.5 0
0
14 Logic Display~
6 694 373 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Z
-4 -22 3 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
44173.5 0
0
14 Logic Display~
6 695 294 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Y
-4 -20 3 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
44173.5 0
0
14 Logic Display~
6 692 206 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 X
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
44173.5 0
0
8 4-In OR~
219 583 391 0 5 22
0 5 4 3 2 9
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
6435 0 0
2
44173.5 0
0
8 4-In OR~
219 581 311 0 5 22
0 6 4 2 2 10
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
5283 0 0
2
44173.5 0
0
8 4-In OR~
219 581 226 0 5 22
0 8 3 7 2 11
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
6874 0 0
2
44173.5 0
0
15
0 4 2 0 0 4096 0 0 12 9 0 2
338 405
566 405
0 3 3 0 0 4224 0 0 12 11 0 3
353 397
566 397
566 396
2 0 4 0 0 4096 0 12 0 0 7 3
566 387
388 387
388 307
1 1 5 0 0 8320 0 7 12 0 0 5
297 243
297 262
537 262
537 378
566 378
4 0 2 0 0 0 0 13 0 0 9 2
564 325
338 325
3 0 2 0 0 0 0 13 0 0 9 3
564 316
564 315
338 315
1 2 4 0 0 8320 0 5 13 0 0 3
299 322
299 307
564 307
1 1 6 0 0 8320 0 6 13 0 0 3
298 285
298 298
564 298
1 4 2 0 0 8320 0 1 14 0 0 4
300 479
338 479
338 240
564 240
1 3 7 0 0 12416 0 2 14 0 0 4
299 436
346 436
346 231
564 231
1 2 3 0 0 0 0 3 14 0 0 4
298 397
353 397
353 222
564 222
1 1 8 0 0 12416 0 4 14 0 0 4
298 359
360 359
360 213
564 213
1 5 9 0 0 4224 0 9 12 0 0 2
694 391
616 391
1 5 10 0 0 8336 0 10 13 0 0 3
695 312
695 311
614 311
1 5 11 0 0 8320 0 11 14 0 0 3
692 224
692 226
614 226
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
