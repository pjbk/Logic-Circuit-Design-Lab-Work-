CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 290 346 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3641 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 281 284 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3104 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 276 219 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3296 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 1062 286 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 1041 97 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
5.89886e-315 0
0
8 4-In OR~
219 1021 304 0 5 22
0 7 6 5 4 2
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3371 0 0
2
5.89886e-315 0
0
8 4-In OR~
219 997 115 0 5 22
0 10 9 8 4 3
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
7311 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 892 401 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 895 345 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3526 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 894 303 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4129 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 892 243 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6278 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 890 196 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 887 158 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8323 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 882 110 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 878 56 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7622 0 0
2
5.89886e-315 0
0
9 Inverter~
13 341 316 0 2 22
0 12 15
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
816 0 0
2
5.89886e-315 0
0
9 Inverter~
13 340 259 0 2 22
0 13 16
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4656 0 0
2
5.89886e-315 0
0
9 Inverter~
13 339 203 0 2 22
0 14 17
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
6356 0 0
2
5.89886e-315 0
0
5 7415~
219 713 423 0 4 22
0 14 13 12 4
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
7479 0 0
2
5.89886e-315 0
0
5 7415~
219 712 373 0 4 22
0 14 13 15 5
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
5690 0 0
2
5.89886e-315 0
0
5 7415~
219 710 324 0 4 22
0 14 16 12 6
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
5617 0 0
2
5.89886e-315 0
0
5 7415~
219 712 274 0 4 22
0 14 16 15 8
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
3903 0 0
2
5.89886e-315 0
0
5 7415~
219 709 224 0 4 22
0 17 13 12 7
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
4452 0 0
2
5.89886e-315 0
0
5 7415~
219 706 175 0 4 22
0 17 13 15 9
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
6282 0 0
2
5.89886e-315 0
0
5 7415~
219 704 127 0 4 22
0 17 16 12 10
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
7187 0 0
2
5.89886e-315 0
0
5 7415~
219 702 78 0 4 22
0 17 16 15 11
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
6866 0 0
2
5.89886e-315 0
0
45
1 5 2 0 0 4224 0 4 6 0 0 2
1062 304
1054 304
1 5 3 0 0 4224 0 5 7 0 0 2
1041 115
1030 115
0 4 4 0 0 8192 0 0 6 11 0 5
858 423
858 329
996 329
996 318
1004 318
0 3 5 0 0 8320 0 0 6 12 0 5
808 373
808 280
991 280
991 309
1004 309
0 2 6 0 0 8320 0 0 6 13 0 5
810 324
810 285
996 285
996 300
1004 300
0 1 7 0 0 8320 0 0 6 15 0 3
792 224
792 291
1004 291
0 4 4 0 0 4224 0 0 7 11 0 5
843 423
843 138
967 138
967 129
980 129
0 3 8 0 0 8192 0 0 7 14 0 5
829 274
829 133
972 133
972 120
980 120
0 2 9 0 0 8320 0 0 7 16 0 5
815 175
815 89
967 89
967 111
980 111
0 1 10 0 0 8320 0 0 7 17 0 5
787 127
787 94
972 94
972 102
980 102
1 4 4 0 0 0 0 8 19 0 0 3
892 419
892 423
734 423
1 4 5 0 0 0 0 9 20 0 0 3
895 363
895 373
733 373
1 4 6 0 0 0 0 10 21 0 0 4
894 321
810 321
810 324
731 324
1 4 8 0 0 8320 0 11 22 0 0 3
892 261
892 274
733 274
1 4 7 0 0 0 0 12 23 0 0 3
890 214
890 224
730 224
1 4 9 0 0 0 0 13 24 0 0 6
887 176
815 176
815 175
726 175
726 175
727 175
1 4 10 0 0 0 0 14 25 0 0 4
882 128
787 128
787 127
725 127
1 4 11 0 0 8336 0 15 26 0 0 5
878 74
878 78
722 78
722 78
723 78
0 3 12 0 0 8192 0 0 19 37 0 3
398 330
398 432
689 432
0 2 13 0 0 8192 0 0 19 35 0 3
419 175
419 423
689 423
0 1 14 0 0 8192 0 0 19 30 0 3
449 274
449 414
689 414
0 3 15 0 0 8192 0 0 20 43 0 3
502 316
502 382
688 382
0 2 13 0 0 0 0 0 20 35 0 3
567 175
567 373
688 373
0 1 14 0 0 0 0 0 20 30 0 3
559 274
559 364
688 364
0 3 12 0 0 0 0 0 21 37 0 3
672 330
672 333
686 333
0 2 16 0 0 4224 0 0 21 44 0 3
581 78
581 324
686 324
0 1 14 0 0 0 0 0 21 30 0 3
577 274
577 315
686 315
0 3 15 0 0 4096 0 0 22 43 0 3
604 87
604 283
688 283
0 2 16 0 0 0 0 0 22 44 0 3
623 78
623 274
688 274
0 1 14 0 0 8320 0 0 22 42 0 5
300 219
300 274
680 274
680 265
688 265
0 3 12 0 0 0 0 0 23 37 0 2
672 233
685 233
0 2 13 0 0 0 0 0 23 35 0 3
609 175
609 224
685 224
0 1 17 0 0 4096 0 0 23 45 0 3
614 69
614 215
685 215
0 3 15 0 0 0 0 0 24 43 0 3
633 87
633 184
682 184
0 2 13 0 0 8320 0 0 24 41 0 3
317 284
317 175
682 175
0 1 17 0 0 0 0 0 24 45 0 3
643 69
643 166
682 166
0 3 12 0 0 4224 0 0 25 40 0 4
318 330
672 330
672 136
680 136
0 2 16 0 0 0 0 0 25 44 0 3
662 78
662 127
680 127
0 1 17 0 0 0 0 0 25 45 0 3
653 69
653 118
680 118
1 1 12 0 0 0 0 1 16 0 0 4
302 346
318 346
318 316
326 316
1 1 13 0 0 0 0 2 17 0 0 4
293 284
317 284
317 259
325 259
1 1 14 0 0 0 0 3 18 0 0 4
288 219
316 219
316 203
324 203
2 3 15 0 0 8320 0 16 26 0 0 4
362 316
512 316
512 87
678 87
2 2 16 0 0 0 0 17 26 0 0 4
361 259
517 259
517 78
678 78
2 1 17 0 0 4224 0 18 26 0 0 4
360 203
522 203
522 69
678 69
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
428 455 665 479
438 463 654 479
27 Full Adder with decoder 3x8
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
