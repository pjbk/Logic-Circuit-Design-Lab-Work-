CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 198 487 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 S1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43653.8 1
0
13 Logic Switch~
5 271 492 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 S0
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43653.8 0
0
13 Logic Switch~
5 124 289 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43653.8 1
0
13 Logic Switch~
5 121 371 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I3
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43653.8 0
0
13 Logic Switch~
5 121 209 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43653.8 0
0
13 Logic Switch~
5 123 127 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43653.8 0
0
9 Inverter~
13 268 432 0 2 22
0 6 8
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
8901 0 0
2
43653.8 0
0
9 Inverter~
13 195 429 0 2 22
0 7 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7361 0 0
2
43653.8 0
0
14 Logic Display~
6 862 170 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43653.8 0
0
5 7415~
219 399 298 0 4 22
0 3 7 8 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
972 0 0
2
43653.8 1
0
5 7415~
219 401 380 0 4 22
0 2 7 6 11
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
3472 0 0
2
43653.8 0
0
5 7415~
219 400 218 0 4 22
0 4 9 6 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
9998 0 0
2
43653.8 0
0
5 7415~
219 398 136 0 4 22
0 5 9 8 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
3536 0 0
2
43653.8 0
0
8 4-In OR~
219 665 216 0 5 22
0 14 13 12 11 10
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
4597 0 0
2
43653.8 0
0
19
1 1 2 0 0 4224 0 11 4 0 0 2
377 371
133 371
1 1 3 0 0 4224 0 10 3 0 0 2
375 289
136 289
1 1 4 0 0 4224 0 12 5 0 0 2
376 209
133 209
1 1 5 0 0 4224 0 13 6 0 0 2
374 127
135 127
3 0 6 0 0 4096 0 11 0 0 10 2
377 389
317 389
2 0 7 0 0 4096 0 11 0 0 8 2
377 380
236 380
3 0 8 0 0 4096 0 10 0 0 13 2
375 307
271 307
0 2 7 0 0 8320 0 0 10 9 0 4
198 456
236 456
236 298
375 298
1 1 7 0 0 0 0 1 8 0 0 3
199 474
198 474
198 447
0 3 6 0 0 8320 0 0 12 11 0 4
271 459
317 459
317 227
376 227
1 1 6 0 0 0 0 2 7 0 0 3
272 479
271 479
271 450
2 0 9 0 0 4096 0 12 0 0 14 2
376 218
198 218
2 3 8 0 0 4224 0 7 13 0 0 3
271 414
271 145
374 145
2 2 9 0 0 4224 0 8 13 0 0 3
198 411
198 136
374 136
1 5 10 0 0 8320 0 9 14 0 0 3
862 188
862 216
698 216
4 4 11 0 0 4224 0 11 14 0 0 4
422 380
635 380
635 230
648 230
4 3 12 0 0 4224 0 10 14 0 0 4
420 298
640 298
640 221
648 221
4 2 13 0 0 4224 0 12 14 0 0 4
421 218
640 218
640 212
648 212
4 1 14 0 0 4224 0 13 14 0 0 4
419 136
640 136
640 203
648 203
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
