CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 81 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 177 457 274
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 101 412 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 bin
-48 -9 -27 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
364 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 107 242 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 y
-39 -12 -32 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3656 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 109 137 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 x
-42 -6 -35 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3131 0 0
2
5.89774e-315 0
0
9 Inverter~
13 668 241 0 2 22
0 8 7
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
6772 0 0
2
5.89774e-315 0
0
9 Inverter~
13 201 335 0 2 22
0 9 10
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9557 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1064 287 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5789 0 0
2
5.89774e-315 0
0
14 Logic Display~
6 1076 142 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7328 0 0
2
5.89774e-315 0
0
8 2-In OR~
219 850 305 0 3 22
0 4 5 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4799 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 765 250 0 3 22
0 7 6 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9196 0 0
2
5.89774e-315 0
0
9 2-In AND~
219 324 326 0 3 22
0 11 10 5
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3857 0 0
2
5.89774e-315 0
0
6 74136~
219 298 147 0 3 22
0 9 11 8
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7125 0 0
2
5.89774e-315 0
0
6 74136~
219 649 160 0 3 22
0 8 6 2
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3641 0 0
2
5.89774e-315 0
0
14
3 1 2 0 0 4224 0 12 7 0 0 2
682 160
1076 160
3 1 3 0 0 4224 0 8 6 0 0 2
883 305
1064 305
3 1 4 0 0 8320 0 9 8 0 0 4
786 250
829 250
829 296
837 296
3 2 5 0 0 4224 0 10 8 0 0 4
345 326
822 326
822 314
837 314
2 0 6 0 0 4096 0 9 0 0 8 2
741 259
625 259
2 1 7 0 0 4224 0 4 9 0 0 2
689 241
741 241
0 1 8 0 0 8192 0 0 4 9 0 3
432 147
432 241
653 241
1 2 6 0 0 4224 0 1 12 0 0 4
113 412
625 412
625 169
633 169
3 1 8 0 0 4224 0 11 12 0 0 4
331 147
625 147
625 151
633 151
0 1 9 0 0 4096 0 0 5 14 0 3
166 137
166 335
186 335
2 2 10 0 0 8320 0 5 10 0 0 2
222 335
300 335
1 0 11 0 0 8192 0 10 0 0 13 4
300 317
289 317
289 242
274 242
1 2 11 0 0 4224 0 2 11 0 0 4
119 242
274 242
274 156
282 156
1 1 9 0 0 4224 0 3 11 0 0 4
121 137
274 137
274 138
282 138
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1026 132 1055 156
1036 140 1044 156
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1005 271 1058 295
1015 279 1047 295
4 bout
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
