CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
14 Logic Display~
6 150 87 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
44174.7 23
0
14 Logic Display~
6 322 85 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
44174.7 22
0
14 Logic Display~
6 472 82 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
44174.7 21
0
14 Logic Display~
6 635 80 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
44174.7 20
0
9 2-In AND~
219 601 356 0 3 22
0 10 23 21
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
754 0 0
2
44174.7 19
0
9 2-In AND~
219 600 420 0 3 22
0 4 22 20
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9767 0 0
2
44174.7 18
0
9 2-In AND~
219 440 437 0 3 22
0 20 5 18
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U5C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7978 0 0
2
44174.7 17
0
9 2-In AND~
219 440 371 0 3 22
0 21 11 19
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U5D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3142 0 0
2
44174.7 16
0
9 2-In AND~
219 290 453 0 3 22
0 18 6 16
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U6A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3284 0 0
2
44174.7 15
0
9 2-In AND~
219 286 386 0 3 22
0 19 9 17
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U6B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
659 0 0
2
44174.7 14
0
9 2-In AND~
219 117 469 0 3 22
0 16 7 33
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U6C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 2 0
1 U
3800 0 0
2
44174.7 13
0
9 2-In AND~
219 115 400 0 3 22
0 17 8 32
0
0 0 608 512
6 74LS08
-21 -24 21 -16
3 U6D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 2 0
1 U
6792 0 0
2
44174.7 12
0
8 2-In OR~
219 697 292 0 3 22
0 23 22 3
0
0 0 608 602
6 74LS32
-21 -24 21 -16
3 U7A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3701 0 0
2
44174.7 11
0
8 2-In OR~
219 524 296 0 3 22
0 21 20 12
0
0 0 608 602
6 74LS32
-21 -24 21 -16
3 U7B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6316 0 0
2
44174.7 10
0
8 2-In OR~
219 363 297 0 3 22
0 19 18 13
0
0 0 608 602
6 74LS32
-21 -24 21 -16
3 U7C
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8734 0 0
2
44174.7 9
0
8 2-In OR~
219 202 313 0 3 22
0 17 16 14
0
0 0 608 602
6 74LS32
-21 -24 21 -16
3 U7D
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7988 0 0
2
44174.7 8
0
9 Inverter~
13 764 250 0 2 22
0 15 2
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U8A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3217 0 0
2
44174.7 7
0
5 4027~
219 698 202 0 7 32
0 30 3 2 3 31 4 10
0
0 0 4704 90
4 4027
7 -60 35 -52
3 U1A
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
3965 0 0
2
44174.7 6
0
5 4027~
219 525 202 0 7 32
0 28 12 2 12 29 5 11
0
0 0 4704 90
4 4027
7 -60 35 -52
3 U1B
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
8239 0 0
2
44174.7 5
0
5 4027~
219 363 207 0 7 32
0 26 13 2 13 27 6 9
0
0 0 4704 90
4 4027
7 -60 35 -52
3 U2A
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
828 0 0
2
44174.7 4
0
5 4027~
219 198 207 0 7 32
0 24 14 2 14 25 7 8
0
0 0 4704 90
4 4027
7 -60 35 -52
3 U2B
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
6187 0 0
2
44174.7 3
0
13 Logic Switch~
5 921 250 0 1 11
0 15
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7107 0 0
2
44174.7 2
0
13 Logic Switch~
5 846 365 0 1 11
0 23
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6433 0 0
2
44174.7 1
0
13 Logic Switch~
5 854 429 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
44174.7 0
0
41
3 0 2 0 0 16 0 18 0 0 18 4
700 203
700 245
683 245
683 250
0 3 3 0 0 16 0 0 13 3 0 2
700 211
700 262
4 2 3 0 0 16 0 18 18 0 0 4
709 203
709 211
691 211
691 203
6 1 4 0 0 16 0 18 6 0 0 5
709 149
709 135
639 135
639 411
620 411
6 2 5 0 0 16 0 19 7 0 0 5
536 149
536 135
479 135
479 446
460 446
6 2 6 0 0 16 0 20 9 0 0 5
374 154
374 140
329 140
329 462
310 462
6 2 7 0 0 16 0 21 11 0 0 5
209 154
209 145
156 145
156 478
137 478
1 0 8 0 0 16 0 1 0 0 9 2
150 105
150 150
7 2 8 0 0 16 0 21 12 0 0 5
191 160
191 150
149 150
149 409
135 409
1 0 9 0 0 16 0 2 0 0 11 4
322 103
322 145
323 145
323 150
7 2 9 0 0 16 0 20 10 0 0 5
356 160
356 150
320 150
320 395
306 395
1 0 10 0 0 16 0 4 0 0 13 4
635 98
635 140
636 140
636 145
7 1 10 0 0 16 0 18 5 0 0 5
691 155
691 145
630 145
630 347
621 347
1 0 11 0 0 16 0 3 0 0 15 4
472 100
472 140
476 140
476 145
7 2 11 0 0 16 0 19 8 0 0 5
518 155
518 145
474 145
474 380
460 380
3 0 2 0 0 16 0 19 0 0 18 2
527 203
527 250
3 0 2 0 0 16 0 20 0 0 18 2
365 208
365 250
3 2 2 0 0 16 0 21 17 0 0 3
200 208
200 250
749 250
0 3 12 0 0 16 0 0 14 20 0 2
527 211
527 266
4 2 12 0 0 16 0 19 19 0 0 4
536 203
536 211
518 211
518 203
0 3 13 0 0 16 0 0 15 22 0 2
366 216
366 267
4 2 13 0 0 16 0 20 20 0 0 4
374 208
374 216
356 216
356 208
4 3 14 0 0 16 0 21 16 0 0 4
209 208
209 277
205 277
205 283
2 3 14 0 0 16 0 21 16 0 0 4
191 208
191 282
205 282
205 283
1 1 15 0 0 16 0 17 22 0 0 2
785 250
907 250
2 0 16 0 0 16 0 16 0 0 28 2
196 329
196 453
1 0 17 0 0 16 0 16 0 0 29 2
214 329
214 386
3 1 16 0 0 16 0 9 11 0 0 4
265 453
146 453
146 460
137 460
3 1 17 0 0 16 0 10 12 0 0 4
261 386
144 386
144 391
135 391
2 0 18 0 0 16 0 15 0 0 32 2
357 313
357 437
1 0 19 0 0 16 0 15 0 0 33 2
375 313
375 371
3 1 18 0 0 16 0 7 9 0 0 4
415 437
319 437
319 444
310 444
3 1 19 0 0 16 0 8 10 0 0 4
415 371
315 371
315 377
306 377
2 0 20 0 0 16 0 14 0 0 36 2
518 312
518 420
1 0 21 0 0 16 0 14 0 0 37 2
536 312
536 356
3 1 20 0 0 16 0 6 7 0 0 4
575 420
469 420
469 428
460 428
3 1 21 0 0 16 0 5 8 0 0 4
576 356
469 356
469 362
460 362
2 0 22 0 0 16 0 13 0 0 40 2
691 308
691 429
1 0 23 0 0 16 0 13 0 0 41 2
709 308
709 365
1 2 22 0 0 16 0 24 6 0 0 2
840 429
620 429
1 2 23 0 0 16 0 23 5 0 0 2
832 365
621 365
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
854 348 1011 372
864 356 1000 372
17 Enable down count
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
867 412 1008 436
877 420 997 436
15 Enable up count
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
