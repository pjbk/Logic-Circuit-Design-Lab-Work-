CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 278 331 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6187 0 0
2
44175.5 0
0
13 Logic Switch~
5 281 284 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7107 0 0
2
44175.5 1
0
13 Logic Switch~
5 276 203 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6433 0 0
2
44175.5 2
0
14 Logic Display~
6 908 398 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8559 0 0
2
44175.5 3
0
14 Logic Display~
6 907 347 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
44175.5 4
0
14 Logic Display~
6 906 306 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5697 0 0
2
44175.5 5
0
14 Logic Display~
6 905 246 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
44175.5 6
0
14 Logic Display~
6 905 201 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
44175.5 7
0
14 Logic Display~
6 903 156 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3795 0 0
2
44175.5 8
0
14 Logic Display~
6 903 103 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
44175.5 9
0
14 Logic Display~
6 900 59 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
44175.5 10
0
9 Inverter~
13 341 316 0 2 22
0 11 14
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
6966 0 0
2
44175.5 11
0
9 Inverter~
13 340 259 0 2 22
0 12 15
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9796 0 0
2
44175.5 12
0
9 Inverter~
13 339 203 0 2 22
0 13 16
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
5952 0 0
2
44175.5 13
0
5 7415~
219 713 423 0 4 22
0 13 12 11 3
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
3649 0 0
2
44175.5 14
0
5 7415~
219 712 373 0 4 22
0 13 12 14 4
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
3716 0 0
2
44175.5 15
0
5 7415~
219 710 324 0 4 22
0 13 15 11 5
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
4797 0 0
2
44175.5 16
0
5 7415~
219 712 274 0 4 22
0 13 15 14 6
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
4681 0 0
2
44175.5 17
0
5 7415~
219 709 224 0 4 22
0 16 12 11 7
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
9730 0 0
2
44175.5 18
0
5 7415~
219 706 175 0 4 22
0 16 12 14 8
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
9874 0 0
2
44175.5 19
0
5 7415~
219 704 127 0 4 22
0 16 15 11 9
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
364 0 0
2
44175.5 20
0
5 7415~
219 702 78 0 4 22
0 16 15 14 10
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
3656 0 0
2
44175.5 21
0
36
0 0 2 0 0 4224 0 0 0 0 0 3
1029 116
1029 115
1030 115
1 4 3 0 0 8320 0 4 15 0 0 3
908 416
908 423
734 423
1 4 4 0 0 8320 0 5 16 0 0 3
907 365
907 373
733 373
1 4 5 0 0 4224 0 6 17 0 0 2
906 324
731 324
1 4 6 0 0 8320 0 7 18 0 0 3
905 264
905 274
733 274
1 4 7 0 0 8320 0 8 19 0 0 3
905 219
905 224
730 224
1 4 8 0 0 4224 0 9 20 0 0 4
903 174
726 174
726 175
727 175
1 4 9 0 0 8320 0 10 21 0 0 3
903 121
903 127
725 127
1 4 10 0 0 8320 0 11 22 0 0 5
900 77
900 78
722 78
722 78
723 78
0 3 11 0 0 8192 0 0 15 28 0 3
398 330
398 432
689 432
0 2 12 0 0 8192 0 0 15 26 0 3
419 175
419 423
689 423
0 1 13 0 0 8192 0 0 15 21 0 3
449 274
449 414
689 414
0 3 14 0 0 8192 0 0 16 34 0 3
502 316
502 382
688 382
0 2 12 0 0 0 0 0 16 26 0 3
567 175
567 373
688 373
0 1 13 0 0 0 0 0 16 21 0 3
559 274
559 364
688 364
0 3 11 0 0 0 0 0 17 28 0 3
672 330
672 333
686 333
0 2 15 0 0 4224 0 0 17 35 0 3
581 78
581 324
686 324
0 1 13 0 0 0 0 0 17 21 0 3
577 274
577 315
686 315
0 3 14 0 0 4096 0 0 18 34 0 3
604 87
604 283
688 283
0 2 15 0 0 0 0 0 18 35 0 3
623 78
623 274
688 274
0 1 13 0 0 8320 0 0 18 33 0 5
300 203
300 274
680 274
680 265
688 265
0 3 11 0 0 0 0 0 19 28 0 2
672 233
685 233
0 2 12 0 0 0 0 0 19 26 0 3
609 175
609 224
685 224
0 1 16 0 0 4096 0 0 19 36 0 3
614 69
614 215
685 215
0 3 14 0 0 0 0 0 20 34 0 3
633 87
633 184
682 184
0 2 12 0 0 8320 0 0 20 32 0 3
317 284
317 175
682 175
0 1 16 0 0 0 0 0 20 36 0 3
643 69
643 166
682 166
0 3 11 0 0 4224 0 0 21 31 0 4
318 330
672 330
672 136
680 136
0 2 15 0 0 0 0 0 21 35 0 3
662 78
662 127
680 127
0 1 16 0 0 0 0 0 21 36 0 3
653 69
653 118
680 118
1 1 11 0 0 0 0 1 12 0 0 4
290 331
318 331
318 316
326 316
1 1 12 0 0 0 0 2 13 0 0 4
293 284
317 284
317 259
325 259
1 1 13 0 0 16 0 3 14 0 0 2
288 203
324 203
2 3 14 0 0 8320 0 12 22 0 0 4
362 316
512 316
512 87
678 87
2 2 15 0 0 0 0 13 22 0 0 4
361 259
517 259
517 78
678 78
2 1 16 0 0 4224 0 14 22 0 0 4
360 203
522 203
522 69
678 69
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
519 458 668 482
529 466 657 482
16 3x8 line decoder
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
