CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 239 226 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-31 -7 -24 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
44173.5 0
0
13 Logic Switch~
5 242 296 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-33 -5 -26 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
44173.5 0
0
13 Logic Switch~
5 243 368 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
44173.5 0
0
5 4023~
219 566 146 0 4 22
0 9 7 10 5
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 2 0
1 U
3108 0 0
2
44173.5 0
0
5 4023~
219 568 214 0 4 22
0 9 6 10 4
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 4 0
1 U
4299 0 0
2
44173.5 0
0
5 4023~
219 570 280 0 4 22
0 8 7 10 3
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 4 0
1 U
9672 0 0
2
44173.5 0
0
5 4023~
219 571 359 0 4 22
0 8 6 10 2
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 4 0
1 U
7876 0 0
2
44173.5 0
0
14 Logic Display~
6 637 341 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
44173.5 0
0
14 Logic Display~
6 634 262 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
44173.5 0
0
14 Logic Display~
6 637 196 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -20 7 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
44173.5 0
0
14 Logic Display~
6 636 128 0 1 2
20 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
44173.5 0
0
5 4049~
219 336 368 0 2 22
0 11 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
7678 0 0
2
44173.5 0
0
5 4049~
219 431 296 0 2 22
0 7 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
961 0 0
2
44173.5 0
0
5 4049~
219 430 226 0 2 22
0 9 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
3178 0 0
2
44173.5 0
0
5 4049~
219 335 296 0 2 22
0 12 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3409 0 0
2
44173.5 0
0
5 4049~
219 332 226 0 2 22
0 13 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
3951 0 0
2
44173.5 0
0
21
4 1 2 0 0 12416 0 7 8 0 0 2
598 359
637 359
4 1 3 0 0 4224 0 6 9 0 0 2
597 280
634 280
4 1 4 0 0 4224 0 5 10 0 0 2
595 214
637 214
4 1 5 0 0 4224 0 4 11 0 0 2
593 146
636 146
0 2 6 0 0 4096 0 0 7 6 0 3
490 294
490 359
547 359
2 2 6 0 0 8320 0 13 5 0 0 4
452 296
490 296
490 214
544 214
0 2 7 0 0 4112 0 0 6 8 0 2
398 280
546 280
0 2 7 0 0 4224 0 0 4 14 0 3
398 296
398 146
542 146
0 1 8 0 0 4096 0 0 6 10 0 2
531 271
546 271
2 1 8 0 0 12416 0 14 7 0 0 5
451 226
451 241
531 241
531 350
547 350
0 1 9 0 0 4224 0 0 5 12 0 2
376 205
544 205
0 1 9 0 0 0 0 0 4 13 0 3
376 226
376 137
542 137
2 1 9 0 0 0 0 16 14 0 0 2
353 226
415 226
2 1 7 0 0 0 0 15 13 0 0 2
356 296
416 296
0 3 10 0 0 8192 0 0 5 18 0 2
513 223
544 223
0 3 10 0 0 4096 0 0 6 18 0 2
513 289
546 289
0 3 10 0 0 4096 0 0 7 18 0 2
513 368
547 368
2 3 10 0 0 8320 0 12 4 0 0 4
357 368
513 368
513 155
542 155
1 1 11 0 0 8320 0 3 12 0 0 2
255 368
321 368
1 1 12 0 0 4224 0 2 15 0 0 2
254 296
320 296
1 1 13 0 0 4224 0 16 1 0 0 2
317 226
251 226
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
185 367 286 391
195 375 275 391
10 Enable pin
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
