CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 831 306 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4292 0 0
2
44174.7 0
0
13 Logic Switch~
5 954 254 0 1 11
0 9
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6118 0 0
2
44174.7 1
0
14 Logic Display~
6 793 70 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44174.7 2
0
14 Logic Display~
6 636 75 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
44174.7 3
0
14 Logic Display~
6 511 71 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
44174.7 4
0
14 Logic Display~
6 395 73 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
44174.7 5
0
5 4049~
219 850 254 0 2 22
0 9 11
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U4A
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
7634 0 0
2
44174.7 6
0
9 2-In AND~
219 323 269 0 3 22
0 8 12 16
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 3 0
1 U
523 0 0
2
44174.7 7
0
9 2-In AND~
219 433 281 0 3 22
0 7 13 12
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6748 0 0
2
44174.7 8
0
9 2-In AND~
219 560 289 0 3 22
0 6 14 13
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6901 0 0
2
44174.7 9
0
9 2-In AND~
219 702 297 0 3 22
0 5 15 14
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
842 0 0
2
44174.7 10
0
5 4027~
219 386 227 0 7 32
0 17 12 11 12 18 8 2
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U2B
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3277 0 0
2
44174.7 11
0
5 4027~
219 500 230 0 7 32
0 19 13 11 13 20 7 10
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U2A
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4212 0 0
2
44174.7 12
0
5 4027~
219 623 228 0 7 32
0 21 14 11 14 22 6 3
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U1B
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4720 0 0
2
44174.7 13
0
5 4027~
219 791 230 0 7 32
0 23 15 11 15 24 5 4
0
0 0 4720 602
4 4027
7 -60 35 -52
3 U1A
31 -52 52 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
5551 0 0
2
44174.7 14
0
28
0 7 2 0 0 4096 0 0 12 9 0 3
395 172
395 180
399 180
0 7 3 0 0 4096 0 0 14 11 0 2
636 167
636 181
0 7 4 0 0 8192 0 0 15 12 0 3
793 171
804 171
804 183
6 1 5 0 0 12416 0 15 11 0 0 5
786 177
786 173
731 173
731 288
722 288
6 1 6 0 0 12416 0 14 10 0 0 5
618 175
618 171
589 171
589 280
580 280
6 1 7 0 0 12416 0 13 9 0 0 5
495 177
495 173
462 173
462 272
453 272
6 1 8 0 0 12416 0 12 8 0 0 5
381 174
381 170
352 170
352 260
343 260
1 1 9 0 0 4224 0 7 2 0 0 2
871 254
942 254
1 0 2 0 0 4224 0 6 0 0 0 3
395 91
395 172
399 172
1 7 10 0 0 4224 0 5 13 0 0 4
511 89
511 173
513 173
513 183
1 0 3 0 0 4224 0 4 0 0 0 2
636 93
636 171
1 0 4 0 0 4224 0 3 0 0 0 3
793 88
793 173
804 173
3 0 11 0 0 4096 0 13 0 0 16 4
504 231
504 249
505 249
505 254
3 0 11 0 0 4096 0 14 0 0 16 2
627 229
627 254
3 0 11 0 0 0 0 15 0 0 16 4
795 231
795 249
796 249
796 254
3 2 11 0 0 8320 0 12 7 0 0 3
390 228
390 254
835 254
4 0 12 0 0 4096 0 12 0 0 19 2
381 228
381 281
2 0 12 0 0 0 0 12 0 0 19 2
399 228
399 281
3 2 12 0 0 4224 0 9 8 0 0 4
408 281
352 281
352 278
343 278
4 0 13 0 0 4096 0 13 0 0 22 2
495 231
495 289
2 0 13 0 0 0 0 13 0 0 22 2
513 231
513 289
3 2 13 0 0 4224 0 10 9 0 0 4
535 289
462 289
462 290
453 290
4 0 14 0 0 4096 0 14 0 0 25 2
618 229
618 297
2 0 14 0 0 0 0 14 0 0 25 2
636 229
636 297
3 2 14 0 0 4224 0 11 10 0 0 4
677 297
589 297
589 298
580 298
4 0 15 0 0 4096 0 15 0 0 28 2
786 231
786 306
2 0 15 0 0 0 0 15 0 0 28 2
804 231
804 306
2 1 15 0 0 4224 0 11 1 0 0 2
722 306
819 306
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
