CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 152 231 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
44175.5 0
0
13 Logic Switch~
5 151 160 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
44175.5 1
0
9 Inverter~
13 568 462 0 2 22
0 7 6
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9968 0 0
2
44175.5 2
0
5 7422~
219 440 455 0 5 22
0 6 4 3 5 2
0
0 0 624 180
6 74LS22
-21 -28 21 -20
3 U5A
-8 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 5 0
1 U
9281 0 0
2
44175.5 3
0
14 Logic Display~
6 964 99 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
44175.5 4
0
6 JK RN~
219 882 231 0 6 22
0 9 7 9 2 11 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
7168 0 0
2
44175.5 5
0
6 JK RN~
219 300 238 0 6 22
0 9 10 9 2 12 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3171 0 0
2
44175.5 6
0
6 JK RN~
219 475 237 0 6 22
0 9 8 9 2 13 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
4139 0 0
2
44175.5 7
0
6 JK RN~
219 672 239 0 6 22
0 9 4 9 2 14 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
6435 0 0
2
44175.5 8
0
14 Logic Display~
6 1064 99 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
44175.5 9
0
14 Logic Display~
6 1031 99 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
44175.5 10
0
14 Logic Display~
6 999 99 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
44175.5 11
0
9 Inverter~
13 564 407 0 2 22
0 8 5
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
34 0 0
2
44175.5 12
0
26
0 4 2 0 0 4096 0 0 8 3 0 2
475 291
475 268
0 4 2 0 0 0 0 0 9 3 0 2
672 291
672 270
0 4 2 0 0 4224 0 0 6 4 0 3
300 291
882 291
882 262
5 4 2 0 0 0 0 4 7 0 0 3
413 455
300 455
300 269
0 3 3 0 0 8320 0 0 4 11 0 5
946 214
946 442
474 442
474 461
464 461
0 2 4 0 0 4224 0 0 4 18 0 3
539 220
539 449
464 449
2 4 5 0 0 4224 0 13 4 0 0 4
549 407
474 407
474 437
464 437
2 1 6 0 0 4224 0 3 4 0 0 4
553 462
474 462
474 473
464 473
0 1 7 0 0 4224 0 0 3 17 0 3
715 222
715 462
589 462
0 1 8 0 0 8320 0 0 13 19 0 7
339 221
339 420
546 420
546 435
594 435
594 407
585 407
6 1 3 0 0 0 0 6 5 0 0 3
906 214
964 214
964 117
3 0 9 0 0 4096 0 6 0 0 13 3
858 232
821 232
821 214
1 0 9 0 0 4096 0 6 0 0 26 4
858 214
706 214
706 163
633 163
0 2 7 0 0 0 0 0 6 17 0 3
735 222
735 223
851 223
0 1 8 0 0 8336 0 0 10 19 0 4
372 221
372 191
1064 191
1064 117
0 1 4 0 0 8320 0 0 11 18 0 4
570 220
570 174
1031 174
1031 117
6 1 7 0 0 12416 0 9 12 0 0 5
696 222
735 222
735 154
999 154
999 117
6 2 4 0 0 0 0 8 9 0 0 4
499 220
628 220
628 231
641 231
6 2 8 0 0 0 0 7 8 0 0 4
324 221
436 221
436 229
444 229
1 2 10 0 0 4224 0 1 7 0 0 4
164 231
261 231
261 230
269 230
3 0 9 0 0 0 0 7 0 0 26 3
276 239
240 239
240 160
1 0 9 0 0 0 0 7 0 0 26 3
276 221
264 221
264 160
3 0 9 0 0 0 0 8 0 0 26 3
451 238
417 238
417 160
1 0 9 0 0 0 0 8 0 0 26 3
451 220
440 220
440 160
3 0 9 0 0 0 0 9 0 0 26 3
648 240
612 240
612 160
1 1 9 0 0 4224 0 2 9 0 0 4
163 160
633 160
633 222
648 222
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
