CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 749 206 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5156 0 0
2
44174.7 0
0
13 Logic Switch~
5 754 240 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3133 0 0
2
44174.7 1
0
13 Logic Switch~
5 595 249 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5523 0 0
2
44174.7 2
0
13 Logic Switch~
5 592 209 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3746 0 0
2
44174.7 3
0
13 Logic Switch~
5 468 201 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5668 0 0
2
44174.7 4
0
13 Logic Switch~
5 478 249 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5368 0 0
2
44174.7 5
0
13 Logic Switch~
5 332 193 0 1 11
0 14
0
0 0 21360 782
2 0V
-6 -22 8 -14
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8293 0 0
2
44174.7 6
0
13 Logic Switch~
5 334 254 0 1 11
0 13
0
0 0 21360 602
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3232 0 0
2
44174.7 7
0
13 Logic Switch~
5 864 221 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6644 0 0
2
44174.7 8
0
5 4027~
219 262 243 0 7 32
0 15 14 5 13 16 6 17
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U3B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
4978 0 0
2
44174.7 9
0
5 4027~
219 410 248 0 7 32
0 18 11 4 10 19 5 20
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U3A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
9207 0 0
2
44174.7 10
0
5 4027~
219 531 249 0 7 32
0 21 8 3 9 22 4 23
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
6998 0 0
2
44174.7 11
0
5 4027~
219 664 248 0 7 32
0 24 12 2 7 25 3 26
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3175 0 0
2
44174.7 12
0
14 Logic Display~
6 614 104 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3378 0 0
2
44174.7 13
0
14 Logic Display~
6 506 103 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
922 0 0
2
44174.7 14
0
14 Logic Display~
6 380 106 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6891 0 0
2
44174.7 15
0
14 Logic Display~
6 233 105 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5407 0 0
2
44174.7 16
0
16
4 1 0 0 0 0 0 10 8 0 0 3
292 225
333 225
333 241
2 1 0 0 0 0 0 10 7 0 0 3
292 207
332 207
332 205
1 3 2 0 0 8336 0 9 13 0 0 2
852 221
694 221
1 0 3 0 0 4224 0 14 0 0 5 2
614 122
614 230
6 3 3 0 0 0 0 13 12 0 0 4
640 230
569 230
569 222
561 222
1 6 4 0 0 4096 0 15 12 0 0 5
506 121
506 188
499 188
499 231
507 231
1 0 5 0 0 4096 0 16 0 0 16 4
380 124
380 187
368 187
368 230
1 6 6 0 0 4224 0 17 10 0 0 3
233 123
233 225
238 225
4 1 7 0 0 4224 0 13 2 0 0 4
694 230
727 230
727 240
742 240
1 2 8 0 0 8320 0 4 12 0 0 4
580 209
567 209
567 213
561 213
4 1 9 0 0 8320 0 12 3 0 0 4
561 231
565 231
565 249
583 249
4 1 10 0 0 8320 0 11 6 0 0 4
440 230
452 230
452 249
466 249
1 2 11 0 0 8320 0 5 11 0 0 4
456 201
448 201
448 212
440 212
1 2 12 0 0 4224 0 1 13 0 0 4
737 206
702 206
702 212
694 212
6 3 4 0 0 4224 0 12 11 0 0 6
507 231
456 231
456 224
448 224
448 221
440 221
6 3 5 0 0 4224 0 11 10 0 0 6
386 230
313 230
313 217
300 217
300 216
292 216
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
