CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 210 190 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 202 263 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 436 98 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
43549.5 0
0
14 Logic Display~
6 567 101 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
43549.5 0
0
14 Logic Display~
6 697 99 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
43549.5 0
0
14 Logic Display~
6 843 95 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89886e-315 0
0
12 D Flip-Flop~
219 769 226 0 4 9
0 4 3 8 7
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8901 0 0
2
5.89886e-315 0
0
12 D Flip-Flop~
219 652 226 0 4 9
0 5 3 9 4
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.89886e-315 0
0
12 D Flip-Flop~
219 511 226 0 4 9
0 6 3 10 5
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89886e-315 0
0
12 D Flip-Flop~
219 388 226 0 4 9
0 2 3 11 6
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
5.89886e-315 0
0
15
1 1 2 0 0 4224 0 1 10 0 0 2
222 190
364 190
2 0 3 0 0 8192 0 10 0 0 5 3
364 208
346 208
346 263
2 0 3 0 0 0 0 8 0 0 5 3
628 208
615 208
615 263
2 0 3 0 0 0 0 9 0 0 5 3
487 208
474 208
474 263
2 1 3 0 0 12416 0 7 2 0 0 4
745 208
686 208
686 263
214 263
1 0 4 0 0 4224 0 5 0 0 13 2
697 117
697 190
1 0 5 0 0 4096 0 4 0 0 14 2
567 119
567 190
1 0 6 0 0 4096 0 3 0 0 15 2
436 116
436 190
1 4 7 0 0 4224 0 6 7 0 0 3
843 113
843 190
793 190
2 0 3 0 0 0 0 10 0 0 0 3
364 208
356 208
356 263
2 0 3 0 0 0 0 9 0 0 0 3
487 208
481 208
481 263
2 0 3 0 0 0 0 8 0 0 0 3
628 208
621 208
621 263
4 1 4 0 0 128 0 8 7 0 0 2
676 190
745 190
4 1 5 0 0 4224 0 9 8 0 0 2
535 190
628 190
4 1 6 0 0 4224 0 10 9 0 0 2
412 190
487 190
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
