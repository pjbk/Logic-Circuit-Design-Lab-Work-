CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 245 271 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43550.5 3
0
13 Logic Switch~
5 246 297 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43550.5 2
0
13 Logic Switch~
5 251 376 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43550.5 1
0
13 Logic Switch~
5 253 403 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43550.5 0
0
13 Logic Switch~
5 248 191 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43550.5 1
0
13 Logic Switch~
5 244 223 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43550.5 0
0
13 Logic Switch~
5 247 122 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
43550.5 0
0
13 Logic Switch~
5 245 95 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7361 0 0
2
43550.5 0
0
14 Logic Display~
6 1001 358 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43550.5 0
0
14 Logic Display~
6 997 279 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43550.5 0
0
14 Logic Display~
6 998 195 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43550.5 0
0
14 Logic Display~
6 998 76 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43550.5 0
0
6 74136~
219 817 388 0 3 22
0 9 8 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3536 0 0
2
43550.5 0
0
6 74136~
219 816 305 0 3 22
0 7 6 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4597 0 0
2
43550.5 0
0
6 74136~
219 815 224 0 3 22
0 4 5 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3835 0 0
2
43550.5 0
0
6 74136~
219 813 125 0 3 22
0 2 3 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3670 0 0
2
43550.5 0
0
9 2-In AND~
219 418 426 0 3 22
0 18 18 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5616 0 0
2
43550.5 0
0
9 2-In AND~
219 422 331 0 3 22
0 20 20 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9323 0 0
2
43550.5 0
0
9 2-In AND~
219 425 247 0 3 22
0 22 22 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
317 0 0
2
43550.5 0
0
9 2-In AND~
219 424 167 0 3 22
0 25 24 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3108 0 0
2
43550.5 0
0
6 74136~
219 415 285 0 3 22
0 20 21 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4299 0 0
2
43550.5 1
0
6 74136~
219 409 382 0 3 22
0 18 19 8
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9672 0 0
2
43550.5 0
0
6 74136~
219 417 211 0 3 22
0 22 23 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7876 0 0
2
43550.5 0
0
6 74136~
219 417 125 0 3 22
0 25 24 2
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6369 0 0
2
43550.5 0
0
6 74S182
133 637 244 0 14 29
0 2 10 4 11 6 12 8 13 3
26 27 5 7 9
0
0 0 4848 0
6 74S182
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 15 14 2 1 4 3 13
7 10 9 11 12 6 5 15 14 2
1 4 3 13 7 10 9 11 12 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
43550.5 0
0
36
1 0 2 0 0 4224 0 16 0 0 9 4
797 116
468 116
468 153
463 153
2 9 3 0 0 4224 0 16 25 0 0 4
797 134
683 134
683 217
669 217
1 0 4 0 0 12416 0 15 0 0 11 5
799 215
679 215
679 197
472 197
472 235
2 12 5 0 0 4224 0 15 25 0 0 4
799 233
683 233
683 262
669 262
2 0 6 0 0 4224 0 14 0 0 13 3
800 314
471 314
471 253
1 13 7 0 0 4224 0 14 25 0 0 4
800 296
683 296
683 271
669 271
2 0 8 0 0 4224 0 13 0 0 15 4
801 397
596 397
596 359
586 359
14 1 9 0 0 4224 0 25 13 0 0 4
669 280
793 280
793 379
801 379
1 3 2 0 0 0 0 25 24 0 0 4
599 217
463 217
463 125
450 125
2 3 10 0 0 4224 0 25 20 0 0 4
599 226
455 226
455 167
445 167
3 3 4 0 0 0 0 25 23 0 0 4
599 235
458 235
458 211
450 211
4 3 11 0 0 4224 0 25 19 0 0 4
599 244
454 244
454 247
446 247
5 3 6 0 0 0 0 25 21 0 0 4
599 253
456 253
456 285
448 285
6 3 12 0 0 4224 0 25 18 0 0 4
599 262
453 262
453 331
443 331
3 7 8 0 0 0 0 22 25 0 0 4
442 382
586 382
586 271
599 271
3 8 13 0 0 4224 0 17 25 0 0 4
439 426
591 426
591 280
599 280
1 3 14 0 0 8320 0 9 13 0 0 3
1001 376
1001 388
850 388
1 3 15 0 0 8320 0 10 14 0 0 3
997 297
997 305
849 305
1 3 16 0 0 8320 0 11 15 0 0 3
998 213
998 224
848 224
1 3 17 0 0 8320 0 12 16 0 0 3
998 94
998 125
846 125
2 0 18 0 0 4096 0 17 0 0 24 3
394 435
319 435
319 373
1 0 18 0 0 0 0 17 0 0 24 3
394 417
376 417
376 373
2 1 19 0 0 4224 0 22 4 0 0 4
393 391
274 391
274 403
265 403
1 1 18 0 0 4224 0 22 3 0 0 4
393 373
272 373
272 376
263 376
2 0 20 0 0 8192 0 18 0 0 28 3
398 340
356 340
356 276
1 0 20 0 0 0 0 18 0 0 28 3
398 322
374 322
374 276
2 1 21 0 0 4224 0 21 2 0 0 4
399 294
267 294
267 297
258 297
1 1 20 0 0 4224 0 21 1 0 0 4
399 276
266 276
266 271
257 271
2 0 22 0 0 4096 0 19 0 0 32 3
401 256
305 256
305 191
1 0 22 0 0 0 0 19 0 0 32 3
401 238
362 238
362 191
1 2 23 0 0 4224 0 6 23 0 0 4
256 223
393 223
393 220
401 220
1 1 22 0 0 4224 0 5 23 0 0 4
260 191
393 191
393 202
401 202
2 0 24 0 0 4096 0 20 0 0 35 3
400 176
310 176
310 122
0 1 25 0 0 4096 0 0 20 36 0 3
353 95
353 158
400 158
1 2 24 0 0 4224 0 7 24 0 0 4
259 122
393 122
393 134
401 134
1 1 25 0 0 4224 0 8 24 0 0 4
257 95
393 95
393 116
401 116
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
