CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 950 343 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 994 230 0 1 11
0 7
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 808 102 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 683 105 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 546 101 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 360 103 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 D3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.89886e-315 0
0
9 2-In AND~
219 497 184 0 3 22
0 8 3 4
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4139 0 0
2
5.89886e-315 0
0
9 Inverter~
13 888 234 0 2 22
0 7 10
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U2A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 0 0
1 U
6435 0 0
2
5.89886e-315 0
0
9 Inverter~
13 757 233 0 2 22
0 6 11
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U2A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 0 0
1 U
5283 0 0
2
5.89886e-315 0
0
9 Inverter~
13 617 230 0 2 22
0 3 12
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U2A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 0 0
1 U
6874 0 0
2
5.89886e-315 0
0
9 Inverter~
13 428 227 0 2 22
0 6 13
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U2A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 0 0
1 U
5305 0 0
2
5.89886e-315 0
0
5 4027~
219 848 261 0 7 32
0 14 2 10 2 15 16 6
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 0 0
1 U
34 0 0
2
5.89886e-315 0
0
5 4027~
219 716 260 0 7 32
0 17 5 11 2 18 19 3
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 0 0
1 U
969 0 0
2
5.89886e-315 0
0
5 4027~
219 573 257 0 7 32
0 20 2 12 2 21 22 8
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 0 0
1 U
8402 0 0
2
5.89886e-315 0
0
5 4027~
219 384 254 0 7 32
0 23 4 13 2 24 5 9
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U1A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3751 0 0
2
5.89886e-315 0
0
22
4 0 2 0 0 8192 0 15 0 0 2 3
414 236
414 295
603 295
4 0 2 0 0 8320 0 14 0 0 6 3
603 239
603 303
951 303
2 4 2 0 0 0 0 14 14 0 0 2
603 221
603 239
4 0 2 0 0 0 0 13 0 0 6 3
746 242
746 274
951 274
4 0 2 0 0 0 0 12 0 0 6 2
878 243
951 243
2 1 2 0 0 16 0 12 1 0 0 3
878 225
951 225
951 330
2 0 3 0 0 4224 0 7 0 0 10 3
517 193
655 193
655 230
3 2 4 0 0 8320 0 7 15 0 0 3
472 184
472 218
414 218
6 2 5 0 0 8320 0 15 13 0 0 5
360 236
360 309
798 309
798 224
746 224
1 0 3 0 0 0 0 10 0 0 15 4
638 230
678 230
678 217
683 217
1 0 6 0 0 8320 0 11 0 0 14 4
449 227
449 277
821 277
821 225
1 0 6 0 0 0 0 9 0 0 14 4
778 233
803 233
803 225
808 225
1 1 7 0 0 4224 0 2 8 0 0 4
982 230
917 230
917 234
909 234
1 7 6 0 0 0 0 3 12 0 0 3
808 120
808 225
830 225
1 7 3 0 0 0 0 4 13 0 0 3
683 123
683 224
698 224
1 0 8 0 0 4224 0 5 0 0 17 4
546 119
546 195
545 195
545 221
7 1 8 0 0 0 0 14 7 0 0 4
555 221
526 221
526 175
517 175
7 1 9 0 0 8320 0 15 6 0 0 3
366 218
360 218
360 121
2 3 10 0 0 4224 0 8 12 0 0 2
873 234
878 234
2 3 11 0 0 4224 0 9 13 0 0 2
742 233
746 233
2 3 12 0 0 4224 0 10 14 0 0 2
602 230
603 230
2 3 13 0 0 4224 0 11 15 0 0 2
413 227
414 227
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
